* ring_oscillator_4

.include nand.cir
.include inverter.cir

.subckt ring_oscillator_4 in out vdd vss
x0 in out s1 vdd vss nand
x1 s1 s2 vdd vss inverter tplv=6.841875037250503e-08 tpwv=2.020069000272714e-07 tnln=6.748500505575265e-08 tnwn=1.2982708631199422e-07 tpotv=1.8238276851064712e-09 tnotv=1.8518385504142827e-09 inverter
x2 s2 s3 vdd vss inverter tplv=6.56682836305218e-08 tpwv=2.2388517487937316e-07 tnln=5.848198414696123e-08 tnwn=1.1941685319388114e-07 tpotv=2.039445601596551e-09 tnotv=2.0386922705583474e-09 inverter
x3 s3 s4 vdd vss inverter tplv=6.866315478738094e-08 tpwv=2.1727806900064508e-07 tnln=6.525389618070123e-08 tnwn=1.2880833551064577e-07 tpotv=1.9956881234397057e-09 tnotv=1.7344872727805138e-09 inverter
x4 s4 s5 vdd vss inverter tplv=6.6943362041987e-08 tpwv=1.9675139883049024e-07 tnln=6.521171296156777e-08 tnwn=1.2365594052102037e-07 tpotv=1.881769414272598e-09 tnotv=1.7592760631561992e-09 inverter
x5 s5 s6 vdd vss inverter tplv=7.190490619890986e-08 tpwv=2.2966438122707396e-07 tnln=6.577997117746744e-08 tnwn=1.22335856023147e-07 tpotv=2.0857262024942684e-09 tnotv=1.917611732446583e-09 inverter
x6 s6 s7 vdd vss inverter tplv=6.924170147817239e-08 tpwv=2.2868705009311262e-07 tnln=6.447638452198923e-08 tnwn=1.1967580182463968e-07 tpotv=2.0202506601005467e-09 tnotv=1.9773698595642156e-09 inverter
x7 s7 s8 vdd vss inverter tplv=6.611094160902692e-08 tpwv=2.214635992024352e-07 tnln=7.250430885867909e-08 tnwn=1.233050539616947e-07 tpotv=2.064881387614514e-09 tnotv=1.8657958051243262e-09 inverter
x8 s8 s9 vdd vss inverter tplv=7.098493396086477e-08 tpwv=2.0709023511762748e-07 tnln=7.216489246212652e-08 tnwn=1.3460415432263613e-07 tpotv=1.690508441478464e-09 tnotv=2.072491228366204e-09 inverter
x9 s9 s10 vdd vss inverter tplv=7.026324432876973e-08 tpwv=1.954825038071752e-07 tnln=6.388977718206469e-08 tnwn=1.2939058296075775e-07 tpotv=2.137164514524811e-09 tnotv=1.9167435170482532e-09 inverter
x10 s10 s11 vdd vss inverter tplv=6.826396987633649e-08 tpwv=2.07149066162826e-07 tnln=6.193489181287204e-08 tnwn=1.2353872617659045e-07 tpotv=1.7902398708485618e-09 tnotv=1.9097302521801175e-09 inverter
x11 s11 s12 vdd vss inverter tplv=6.08769924374385e-08 tpwv=2.169981876895304e-07 tnln=7.046388117951652e-08 tnwn=1.1945255482606354e-07 tpotv=1.903301959675877e-09 tnotv=1.827211959019071e-09 inverter
x12 s12 out vdd vss inverter tplv=6.814632701587573e-08 tpwv=2.226318391720804e-07 tnln=6.721370948740749e-08 tnwn=1.3172673110860993e-07 tpotv=1.9314601363845115e-09 tnotv=1.90430984081905e-09 inverter
.ends ring_oscillator_4