*nand

.subckt nand A B out vdd vss
M1 vdd A out vdd tp L=65n W=130n, AS=75.3f AD=75.3f PS=1.23u PD=1.23u
M2 vdd B out vdd tp L=65n W=130n, AS=75.3f AD=75.3f PS=1.23u PD=1.23u
M3 out A C vss tn L=65n W=130n AS=75.3f AD=75.3f PS=1.12u PD=1.23u
M4 C B vss vss tn L=65n W=130n AS=75.3f AD=75.3f PS=1.12u PD=1.23u

*BSIM 4.8.2 models
.model tp pmos level=54 version=4.8.2 toxe=1.95n
.model tn nmos level=54 version=4.8.2 toxe=1.85n

.ends nand
