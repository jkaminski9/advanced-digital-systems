* ring_oscillator_3

.include nand.cir
.include inverter.cir

.subckt ring_oscillator_3 in out vdd vss
x0 in out s1 vdd vss nand
x1 s1 s2 vdd vss inverter tplv=6.360423176896149e-08 tpwv=2.261185467753263e-07 tnln=6.313176400076248e-08 tnwn=1.2563784957597469e-07 tpotv=1.9699559037816043e-09 tnotv=1.7961512641920013e-09 inverter
x2 s2 s3 vdd vss inverter tplv=6.434530485429757e-08 tpwv=1.9284616273439094e-07 tnln=6.613737543025526e-08 tnwn=1.4107157247248497e-07 tpotv=1.942810496398608e-09 tnotv=1.876138492580283e-09 inverter
x3 s3 s4 vdd vss inverter tplv=6.400001701566087e-08 tpwv=1.958114831725454e-07 tnln=6.133098008372927e-08 tnwn=1.2205589356483953e-07 tpotv=1.9446570306771826e-09 tnotv=1.7024821525319392e-09 inverter
x4 s4 s5 vdd vss inverter tplv=7.009547186141391e-08 tpwv=2.1405709198215104e-07 tnln=6.73437285075257e-08 tnwn=1.2877331727277939e-07 tpotv=1.8495323911979724e-09 tnotv=1.7672785219001006e-09 inverter
x5 s5 s6 vdd vss inverter tplv=6.38151024624108e-08 tpwv=2.3265318257880044e-07 tnln=6.537494902202634e-08 tnwn=1.236792406205536e-07 tpotv=2.0077497491547717e-09 tnotv=1.9870991931883824e-09 inverter
x6 s6 s7 vdd vss inverter tplv=6.638188937027301e-08 tpwv=2.3531168929998767e-07 tnln=6.254725255587579e-08 tnwn=1.2603978021983849e-07 tpotv=2.05049057924358e-09 tnotv=1.7354322759459645e-09 inverter
x7 s7 s8 vdd vss inverter tplv=5.831848160274653e-08 tpwv=2.186485767612941e-07 tnln=6.917118039618886e-08 tnwn=1.303896234076744e-07 tpotv=1.82762809584095e-09 tnotv=1.887401190838627e-09 inverter
x8 s8 s9 vdd vss inverter tplv=6.974775730957882e-08 tpwv=2.184150909816076e-07 tnln=6.024258559633635e-08 tnwn=1.3613157114384205e-07 tpotv=1.9648714576066372e-09 tnotv=1.8022901709756305e-09 inverter
x9 s9 s10 vdd vss inverter tplv=6.711873531924019e-08 tpwv=1.9717557518720141e-07 tnln=6.04929162933126e-08 tnwn=1.15853081725485e-07 tpotv=2.0339033472667616e-09 tnotv=1.8931891019329865e-09 inverter
x10 s10 s11 vdd vss inverter tplv=6.225046656230556e-08 tpwv=2.0490505013918172e-07 tnln=6.565447200528881e-08 tnwn=1.3764484189811983e-07 tpotv=1.9634767179986127e-09 tnotv=1.8048157094931152e-09 inverter
x11 s11 s12 vdd vss inverter tplv=6.022635214071597e-08 tpwv=2.1516239397892368e-07 tnln=6.924778856873467e-08 tnwn=1.371385018320087e-07 tpotv=1.8731964745172775e-09 tnotv=1.7342282491598707e-09 inverter
x12 s12 out vdd vss inverter tplv=6.66333709425412e-08 tpwv=2.0496724317315433e-07 tnln=6.935356879920805e-08 tnwn=1.4459106671399878e-07 tpotv=2.0112296842745176e-09 tnotv=1.97132260472238e-09 inverter
.ends ring_oscillator_3