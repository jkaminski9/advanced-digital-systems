* ring_oscillator_7

.include nand.cir
.include inverter.cir

.subckt ring_oscillator_7 in out vdd vss
x0 in out s1 vdd vss nand
x1 s1 s2 vdd vss inverter tplv=6.347162204639886e-08 tpwv=2.1705511765979378e-07 tnln=6.063996409814888e-08 tnwn=1.2705280153492678e-07 tpotv=1.9418529162408575e-09 tnotv=1.879028791402148e-09 inverter
x2 s2 s3 vdd vss inverter tplv=6.950461913060987e-08 tpwv=2.1383702294157324e-07 tnln=7.099569770472933e-08 tnwn=1.2564843684235132e-07 tpotv=1.9518158871937564e-09 tnotv=1.889622590945913e-09 inverter
x3 s3 s4 vdd vss inverter tplv=5.927078584928287e-08 tpwv=2.167921578567536e-07 tnln=6.510377166595967e-08 tnwn=1.1327864224692231e-07 tpotv=1.8750692736627587e-09 tnotv=1.7931815324791376e-09 inverter
x4 s4 s5 vdd vss inverter tplv=5.366443887611063e-08 tpwv=2.1852708402666462e-07 tnln=6.111841310877581e-08 tnwn=1.3341477120733775e-07 tpotv=1.7012742205466864e-09 tnotv=1.8405251936247029e-09 inverter
x5 s5 s6 vdd vss inverter tplv=6.362751773605652e-08 tpwv=2.084143609760649e-07 tnln=6.207084805466726e-08 tnwn=1.3242372974287642e-07 tpotv=1.8554955716571513e-09 tnotv=1.9818764385117594e-09 inverter
x6 s6 s7 vdd vss inverter tplv=6.313088597854042e-08 tpwv=2.0016185943477111e-07 tnln=6.474358112675406e-08 tnwn=1.3391740892644916e-07 tpotv=1.7729883385403936e-09 tnotv=1.8557321203238622e-09 inverter
x7 s7 s8 vdd vss inverter tplv=6.048781995134467e-08 tpwv=2.0790907804561866e-07 tnln=7.062820884496091e-08 tnwn=1.2507841525293656e-07 tpotv=2.107001650579151e-09 tnotv=1.9696126165569325e-09 inverter
x8 s8 s9 vdd vss inverter tplv=6.473930766204344e-08 tpwv=2.1974130851835114e-07 tnln=6.608977350828258e-08 tnwn=1.3104097274564598e-07 tpotv=2.0273524656215437e-09 tnotv=1.878806196074034e-09 inverter
x9 s9 s10 vdd vss inverter tplv=7.087698728367057e-08 tpwv=1.977568409821107e-07 tnln=6.438867517984322e-08 tnwn=1.2661753511844645e-07 tpotv=1.930260877174845e-09 tnotv=1.5915699520012867e-09 inverter
x10 s10 s11 vdd vss inverter tplv=6.588873327711153e-08 tpwv=1.993104914236192e-07 tnln=6.10317820706972e-08 tnwn=1.346495667138438e-07 tpotv=1.7393793987253606e-09 tnotv=1.6501293073920614e-09 inverter
x11 s11 s12 vdd vss inverter tplv=6.612167461661709e-08 tpwv=2.404413530448754e-07 tnln=6.149112259034681e-08 tnwn=1.332266041407413e-07 tpotv=1.953605917600314e-09 tnotv=1.8566095968010175e-09 inverter
x12 s12 out vdd vss inverter tplv=6.05356909104102e-08 tpwv=2.3965680635015963e-07 tnln=6.157264935390164e-08 tnwn=1.2020637195269587e-07 tpotv=1.938983368820938e-09 tnotv=1.8328020472001681e-09 inverter
.ends ring_oscillator_7