* ring_oscillator_0

.include nand.cir
.include inverter.cir

.subckt ring_oscillator_0 in out vdd vss
x0 in out s1 vdd vss nand
x1 s1 s2 vdd vss inverter tplv=6.23522003053471e-08 tpwv=2.1146846558977913e-07 tnln=6.704814621764928e-08 tnwn=1.262798691395377e-07 tpotv=1.837851234118949e-09 tnotv=1.7914121674189902e-09 inverter
x2 s2 s3 vdd vss inverter tplv=6.476872161992865e-08 tpwv=2.3505738122048028e-07 tnln=6.470621021199193e-08 tnwn=1.2962342752235734e-07 tpotv=1.7858009515719441e-09 tnotv=1.6708573296716168e-09 inverter
x3 s3 s4 vdd vss inverter tplv=6.705833127323844e-08 tpwv=2.1306050034429763e-07 tnln=6.194789668591942e-08 tnwn=1.456978385931944e-07 tpotv=2.0328564180616604e-09 tnotv=1.8385856657047455e-09 inverter
x4 s4 s5 vdd vss inverter tplv=7.15576415887617e-08 tpwv=2.231586303358449e-07 tnln=6.110477289041955e-08 tnwn=1.3276767082303066e-07 tpotv=1.975694720358198e-09 tnotv=1.8466099352091424e-09 inverter
x5 s5 s6 vdd vss inverter tplv=6.52402427853921e-08 tpwv=2.0413261509421749e-07 tnln=6.024879871520764e-08 tnwn=1.302742859935055e-07 tpotv=1.8909511927908355e-09 tnotv=1.9252565071492097e-09 inverter
x6 s6 s7 vdd vss inverter tplv=7.341610595353034e-08 tpwv=2.2492376630446666e-07 tnln=6.674243102418105e-08 tnwn=1.2452431353884695e-07 tpotv=1.8680979867255986e-09 tnotv=1.8616009747592118e-09 inverter
x7 s7 s8 vdd vss inverter tplv=6.278421985193326e-08 tpwv=1.929500826861315e-07 tnln=6.866592217536874e-08 tnwn=1.29386969760784e-07 tpotv=1.906890896575531e-09 tnotv=1.8528019267870748e-09 inverter
x8 s8 s9 vdd vss inverter tplv=6.295089766122872e-08 tpwv=2.1304571860628223e-07 tnln=6.64691288018254e-08 tnwn=1.3273038419397323e-07 tpotv=1.87258357069638e-09 tnotv=1.9406329138702376e-09 inverter
x9 s9 s10 vdd vss inverter tplv=5.972005299268035e-08 tpwv=2.1203795815090182e-07 tnln=6.41689035427191e-08 tnwn=1.274276263934543e-07 tpotv=1.841631066734171e-09 tnotv=1.7845637009938222e-09 inverter
x10 s10 s11 vdd vss inverter tplv=6.764113390224009e-08 tpwv=1.9257788614938813e-07 tnln=6.257748477568314e-08 tnwn=1.2866568685198202e-07 tpotv=1.7497291443002814e-09 tnotv=1.8291424203111584e-09 inverter
x11 s11 s12 vdd vss inverter tplv=6.539775106035896e-08 tpwv=1.9797486853220678e-07 tnln=6.4576148513191e-08 tnwn=1.1489497772979768e-07 tpotv=1.948876442496291e-09 tnotv=1.9249155041572785e-09 inverter
x12 s12 out vdd vss inverter tplv=6.704235760115531e-08 tpwv=2.3498722108103203e-07 tnln=6.302595357561696e-08 tnwn=1.3912194954177008e-07 tpotv=2.0698780913402496e-09 tnotv=1.711279337298563e-09 inverter
.ends ring_oscillator_0