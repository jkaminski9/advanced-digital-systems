* run_oscillators

.include ring_oscillator_0.cir
.include ring_oscillator_0.cir
.include ring_oscillator_0.cir
.include ring_oscillator_0.cir
.include ring_oscillator_0.cir
.include ring_oscillator_0.cir
.include ring_oscillator_0.cir
.include ring_oscillator_0.cir

x0 en out0 vdd vss ring_oscillator_0
x1 en out1 vdd vss ring_oscillator_0
x2 en out2 vdd vss ring_oscillator_0
x3 en out3 vdd vss ring_oscillator_0
x4 en out4 vdd vss ring_oscillator_0
x5 en out5 vdd vss ring_oscillator_0
x6 en out6 vdd vss ring_oscillator_0
x7 en out7 vdd vss ring_oscillator_0

*set the temperature
.options temp=40

* supply
V0 vdd vss dc 1.2
V1 vss 0 0
* voltage on the input
Vin0 en 0 pulse(1.2 0 1ns 1ns 20ns 480ns)
.control
tran 0.1n 1000n 0

plot en out0 out1 out2 out3 out4 out5 out6 out7 
.endc
.end
