
module clock_mgmt (
	inclk,
	outclk);	

	input		inclk;
	output		outclk;
endmodule
