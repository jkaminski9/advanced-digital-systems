* ring_oscillator_1

.include nand.cir
.include inverter.cir

.subckt ring_oscillator_1 in out vdd vss
x0 in out s1 vdd vss nand
x1 s1 s2 vdd vss inverter tplv=7.149748928557432e-08 tpwv=2.1830971077358787e-07 tnln=6.923627275891937e-08 tnwn=1.2572009798339532e-07 tpotv=2.0109506224215115e-09 tnotv=1.6887261695287032e-09 inverter
x2 s2 s3 vdd vss inverter tplv=6.307036435888065e-08 tpwv=2.1166651844537173e-07 tnln=6.873541746310734e-08 tnwn=1.3253258436202123e-07 tpotv=1.959152074456548e-09 tnotv=1.7614580932475268e-09 inverter
x3 s3 s4 vdd vss inverter tplv=6.378016660119194e-08 tpwv=2.1394595479982986e-07 tnln=6.547428703328195e-08 tnwn=1.1698340276129675e-07 tpotv=2.0836565188172724e-09 tnotv=1.8329725075363045e-09 inverter
x4 s4 s5 vdd vss inverter tplv=7.47248991713666e-08 tpwv=2.4469471017059804e-07 tnln=6.771662588392048e-08 tnwn=1.4319473324062842e-07 tpotv=1.9447072573083566e-09 tnotv=1.8343995637439298e-09 inverter
x5 s5 s6 vdd vss inverter tplv=6.788826235899495e-08 tpwv=2.1631587063610183e-07 tnln=6.715736526369517e-08 tnwn=1.1623985264140907e-07 tpotv=1.948184862300254e-09 tnotv=1.976974333871644e-09 inverter
x6 s6 s7 vdd vss inverter tplv=6.448618207230565e-08 tpwv=2.0800323633863744e-07 tnln=6.788059530924404e-08 tnwn=1.3230924775992926e-07 tpotv=1.907070383796107e-09 tnotv=1.8833866063598487e-09 inverter
x7 s7 s8 vdd vss inverter tplv=6.725846703243173e-08 tpwv=2.2575692128178362e-07 tnln=5.920231183477416e-08 tnwn=1.3916260411378054e-07 tpotv=1.9461504870035658e-09 tnotv=1.75126835325905e-09 inverter
x8 s8 s9 vdd vss inverter tplv=6.97325766220999e-08 tpwv=2.226248725072245e-07 tnln=6.324440977660698e-08 tnwn=1.3666240072320274e-07 tpotv=2.104910801420505e-09 tnotv=1.8489488373767833e-09 inverter
x9 s9 s10 vdd vss inverter tplv=6.33759141416671e-08 tpwv=2.2110580342920837e-07 tnln=6.631287052591256e-08 tnwn=1.1388390244121873e-07 tpotv=1.940283906446904e-09 tnotv=1.8220360266901891e-09 inverter
x10 s10 s11 vdd vss inverter tplv=6.395378813203456e-08 tpwv=2.214927129823025e-07 tnln=6.762950000182257e-08 tnwn=1.231211129838119e-07 tpotv=1.7408832196998244e-09 tnotv=1.981755761329007e-09 inverter
x11 s11 s12 vdd vss inverter tplv=6.68308830681089e-08 tpwv=2.2013839611520465e-07 tnln=5.956191020357183e-08 tnwn=1.1564781805403405e-07 tpotv=1.9571628587557833e-09 tnotv=1.7915632709237126e-09 inverter
x12 s12 out vdd vss inverter tplv=6.218565390646224e-08 tpwv=2.1213632463928546e-07 tnln=6.300461988778641e-08 tnwn=1.32680418113724e-07 tpotv=1.8947570167652946e-09 tnotv=1.7751503006311021e-09 inverter
.ends ring_oscillator_1