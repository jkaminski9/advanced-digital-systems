* ring_oscillator_6

.include nand.cir
.include inverter.cir

.subckt ring_oscillator_6 in out vdd vss
x0 in out s1 vdd vss nand
x1 s1 s2 vdd vss inverter tplv=6.676584255503658e-08 tpwv=2.1747930315973903e-07 tnln=5.976168071499338e-08 tnwn=1.315196307768361e-07 tpotv=2.018795790726574e-09 tnotv=1.8254052038786258e-09 inverter
x2 s2 s3 vdd vss inverter tplv=6.082786440968002e-08 tpwv=2.0352795293888502e-07 tnln=6.68010486217516e-08 tnwn=1.2906712799333418e-07 tpotv=2.0660631826200035e-09 tnotv=1.866564346323933e-09 inverter
x3 s3 s4 vdd vss inverter tplv=6.11674737252951e-08 tpwv=2.1389919937963411e-07 tnln=6.133751085236636e-08 tnwn=1.3544988585877464e-07 tpotv=1.943418833497238e-09 tnotv=1.8262461214586973e-09 inverter
x4 s4 s5 vdd vss inverter tplv=6.778460559887693e-08 tpwv=2.20916075516665e-07 tnln=7.002193156336077e-08 tnwn=1.2908396238962778e-07 tpotv=1.9286860225944288e-09 tnotv=1.7534592216612737e-09 inverter
x5 s5 s6 vdd vss inverter tplv=6.670432216155773e-08 tpwv=2.3045807817752363e-07 tnln=6.73340513746427e-08 tnwn=1.243661423219843e-07 tpotv=1.9374107681464836e-09 tnotv=1.738906493382605e-09 inverter
x6 s6 s7 vdd vss inverter tplv=6.772577725121437e-08 tpwv=1.9116919282920308e-07 tnln=6.694430211563849e-08 tnwn=1.4306935734096424e-07 tpotv=1.978053802135313e-09 tnotv=1.6727743139222607e-09 inverter
x7 s7 s8 vdd vss inverter tplv=6.307532908465213e-08 tpwv=2.1432380239039664e-07 tnln=5.8075237958803876e-08 tnwn=1.3150105861892968e-07 tpotv=1.9571528851693867e-09 tnotv=1.6535922327594564e-09 inverter
x8 s8 s9 vdd vss inverter tplv=7.080460233504652e-08 tpwv=2.036924546068454e-07 tnln=6.298481664086947e-08 tnwn=1.2602168816763854e-07 tpotv=1.9072000769162328e-09 tnotv=1.7492893475448598e-09 inverter
x9 s9 s10 vdd vss inverter tplv=6.102883989782112e-08 tpwv=2.2553783508464244e-07 tnln=6.300739251412117e-08 tnwn=1.3676577515137103e-07 tpotv=1.9423867046829926e-09 tnotv=1.8091092242154766e-09 inverter
x10 s10 s11 vdd vss inverter tplv=5.892633945165566e-08 tpwv=2.1253381342084382e-07 tnln=6.499813587893636e-08 tnwn=1.3147776874461696e-07 tpotv=2.059342106916543e-09 tnotv=1.8176667073039874e-09 inverter
x11 s11 s12 vdd vss inverter tplv=6.252705553731652e-08 tpwv=2.0226847119483405e-07 tnln=6.489761835171162e-08 tnwn=1.4271378565296963e-07 tpotv=1.7993413099351143e-09 tnotv=1.809702755753779e-09 inverter
x12 s12 out vdd vss inverter tplv=6.485421824005369e-08 tpwv=2.2964892920651585e-07 tnln=6.842565655005192e-08 tnwn=1.0996095835927949e-07 tpotv=2.033011222482332e-09 tnotv=1.7238635244588094e-09 inverter
.ends ring_oscillator_6