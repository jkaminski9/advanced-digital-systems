* ring_oscillator_5

.include nand.cir
.include inverter.cir

.subckt ring_oscillator_5 in out vdd vss
x0 in out s1 vdd vss nand
x1 s1 s2 vdd vss inverter tplv=6.091091675878118e-08 tpwv=2.4239087295970345e-07 tnln=6.594787335267214e-08 tnwn=1.3042132300539929e-07 tpotv=1.8900149158328566e-09 tnotv=1.7371162637526103e-09 inverter
x2 s2 s3 vdd vss inverter tplv=5.778589855948224e-08 tpwv=2.4140284350754317e-07 tnln=6.486720387260334e-08 tnwn=1.4173107152922304e-07 tpotv=1.971513529435067e-09 tnotv=1.8193759197611688e-09 inverter
x3 s3 s4 vdd vss inverter tplv=6.177856046790839e-08 tpwv=1.7048153659298356e-07 tnln=5.937774107028977e-08 tnwn=1.275728291125809e-07 tpotv=2.054937752526971e-09 tnotv=1.908810568986991e-09 inverter
x4 s4 s5 vdd vss inverter tplv=6.824617260969172e-08 tpwv=1.9944754520637057e-07 tnln=6.166676783600938e-08 tnwn=1.2944535592494827e-07 tpotv=1.88113082977022e-09 tnotv=1.8891083811939952e-09 inverter
x5 s5 s6 vdd vss inverter tplv=6.680264817945507e-08 tpwv=2.0592788762950825e-07 tnln=6.825576331493836e-08 tnwn=1.2942062794309758e-07 tpotv=1.9193599584510023e-09 tnotv=1.7605057980397561e-09 inverter
x6 s6 s7 vdd vss inverter tplv=6.926692868780248e-08 tpwv=1.9914482960498552e-07 tnln=6.356526541023442e-08 tnwn=1.2872326713547667e-07 tpotv=2.024707380901796e-09 tnotv=1.685812279217732e-09 inverter
x7 s7 s8 vdd vss inverter tplv=6.484526826124765e-08 tpwv=2.1505637385492763e-07 tnln=6.926669963159388e-08 tnwn=1.3895615986197065e-07 tpotv=1.878566415140211e-09 tnotv=1.8859816648131267e-09 inverter
x8 s8 s9 vdd vss inverter tplv=5.999126756644391e-08 tpwv=2.1656297600987516e-07 tnln=6.476870513107295e-08 tnwn=1.2446551084073957e-07 tpotv=1.821742198724927e-09 tnotv=1.826383573050555e-09 inverter
x9 s9 s10 vdd vss inverter tplv=5.7388739893309446e-08 tpwv=2.1644021454826956e-07 tnln=6.716220633502635e-08 tnwn=1.3022148733799982e-07 tpotv=1.8702283270316825e-09 tnotv=2.0473484156606725e-09 inverter
x10 s10 s11 vdd vss inverter tplv=6.919352519999038e-08 tpwv=2.0311150784041062e-07 tnln=6.577384016191943e-08 tnwn=1.2553761998188326e-07 tpotv=2.0124485636663538e-09 tnotv=2.0553907289328427e-09 inverter
x11 s11 s12 vdd vss inverter tplv=6.737499143878837e-08 tpwv=1.9937437453222855e-07 tnln=6.970542664975073e-08 tnwn=1.25065334969685e-07 tpotv=1.9628848071375157e-09 tnotv=1.762561375360032e-09 inverter
x12 s12 out vdd vss inverter tplv=6.636827047375068e-08 tpwv=2.122884361255234e-07 tnln=7.107403206231412e-08 tnwn=1.3831441815312742e-07 tpotv=1.9592600929995003e-09 tnotv=1.700554656257735e-09 inverter
.ends ring_oscillator_5