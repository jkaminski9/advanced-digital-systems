library ieee;
use ieee.std_logic_1164.all;
use ieee.math_real.all;
use ieee.numeric_std.all;

library ads;
use ads.ads_fixed.all;
use ads.ads_complex_pkg.all;

library vga;
use vga.vga_pkg.all;
use vga.vga_data.all;

package mandlebrot_pkg is
	
	-- Constants and types -- 
	
	constant max_iterations     : integer    := 25;
	constant memory_size        : natural    := natural(log2(real(max_iterations)));
	constant threshold          : ads_sfixed := to_ads_sfixed(4);		
	constant vga_width          : natural    := 1920;
	constant vga_height         : natural    := 1080;
	constant mandlebrot_vga_res : vga_timing := vga_res_default;
	
	constant mandlebrot_xmax    : integer := 3;
	constant mandlebrot_xmin    : integer := -3;
	
	constant mandlebrot_xmax_sfixed    : ads_sfixed := to_ads_sfixed(mandlebrot_xmax);
	constant mandlebrot_xmin_sfixed    : ads_sfixed := to_ads_sfixed(mandlebrot_xmin);

	constant mandlebrot_ymax    : integer := 2;
	constant mandlebrot_ymin    : integer := -2;
	
	constant mandlebrot_ymax_sfixed    : ads_sfixed := to_ads_sfixed(mandlebrot_ymax);
	constant mandlebrot_ymin_sfixed    : ads_sfixed := to_ads_sfixed(mandlebrot_ymin);
		
	constant mandlebrot_delta_x : ads_sfixed := to_ads_sfixed(0.003125); --"00000000000000000011001100110"; -- 4 / 640 = 0.00625
	constant mandlebrot_delta_y : ads_sfixed := to_ads_sfixed(0.003704); -- 4 / 480 = 0.00833

	constant num_pixels     : natural    := vga_height * vga_height;
		
	type map_array is array (0 to max_iterations -1 ) of 
							natural range 0 to 15;					
	
	constant cmap_blue : map_array := (
								15,
								15,
								15,
								15,
								15,
								15,
								15,
								15,
								15,
								15,
								15,
								15,
								15,
								15,
								15,
								15,
								13,
								11,
								9,
								7,
								5,
								3,
								1,
								0,
								0);
								
	constant cmap_red : map_array := (
								0,
								1,
								2,
								3,
								4,
								5,
								6,
								7,
								8,
								9,
								10,
								11,
								12,
								13,
								14,
								15,
								15,
								15,
								15,
								15,
								15,
								15,
								15,
								15,
								0);
	constant cmap_green : map_array := (
								0,
								1,
								2,
								3,
								4,
								5,
								6,
								7,
								8,
								9,
								10,
								11,
								12,
								13,
								14,
								15,
								15,
								15,
								15,
								15,
								15,
								15,
								15,
								15,
								0);	
	type stage_type is
	record
		z: ads_complex;
		c: ads_complex;
		stage_data: natural;
		stage_overflow: boolean;
		stage_valid : boolean;
	end record stage_type;
	
	component edge_detector is
			port (
				signal_in:	in	std_logic;
				clock:		in	std_logic;
				reset:		in	std_logic;
				edge_out:	out	std_logic
			);
		end component edge_detector;
		component seed_fsm is
			port (
				clock:		in	std_logic;
				reset:			in	std_logic;
				toggle:        in std_logic;
				seed :			out	ads_complex
			);
		end component seed_fsm;
		component pipeline_stage is
			generic(
				threshold : ads_sfixed := to_ads_sfixed(4);
				stage_number : natural := 0
			);
			port(
				clock : in std_logic;
				reset : in std_logic;
				enable : in std_logic;
				stage_input : in stage_type;
				stage_output : out stage_type
			);
		end component pipeline_stage;
		
		component pipeline is 
			generic (
				num_stages : positive := 23
			);
			port (
					-- Inputs --
					reset : in std_logic;
					clock : in std_logic;
					enable : in std_logic;
					seed  : in ads_complex;
					z0    : in ads_complex;
					-- Outputs --
					iteration : out natural range 0 to num_stages-1;
					output_valid : out std_logic
			);
		end component pipeline;
	
	type seed_array is array(0 to 1099) of ads_complex;
	
	constant julia_seeds : seed_array := (
(re => to_ads_sfixed(-0.16) , im => to_ads_sfixed(1.0405)),
(re => to_ads_sfixed(-0.16562) , im => to_ads_sfixed(1.032555)),
(re => to_ads_sfixed(-0.17124) , im => to_ads_sfixed(1.02461)),
(re => to_ads_sfixed(-0.17686) , im => to_ads_sfixed(1.016665)),
(re => to_ads_sfixed(-0.18248) , im => to_ads_sfixed(1.00872)),
(re => to_ads_sfixed(-0.1881) , im => to_ads_sfixed(1.000775)),
(re => to_ads_sfixed(-0.19372) , im => to_ads_sfixed(0.99283)),
(re => to_ads_sfixed(-0.19934) , im => to_ads_sfixed(0.984885)),
(re => to_ads_sfixed(-0.20496) , im => to_ads_sfixed(0.97694)),
(re => to_ads_sfixed(-0.21058) , im => to_ads_sfixed(0.968995)),
(re => to_ads_sfixed(-0.2162) , im => to_ads_sfixed(0.96105)),
(re => to_ads_sfixed(-0.22182) , im => to_ads_sfixed(0.953105)),
(re => to_ads_sfixed(-0.22744) , im => to_ads_sfixed(0.94516)),
(re => to_ads_sfixed(-0.23306) , im => to_ads_sfixed(0.937215)),
(re => to_ads_sfixed(-0.23868) , im => to_ads_sfixed(0.92927)),
(re => to_ads_sfixed(-0.2443) , im => to_ads_sfixed(0.921325)),
(re => to_ads_sfixed(-0.24992) , im => to_ads_sfixed(0.91338)),
(re => to_ads_sfixed(-0.25554) , im => to_ads_sfixed(0.905435)),
(re => to_ads_sfixed(-0.26116) , im => to_ads_sfixed(0.89749)),
(re => to_ads_sfixed(-0.26678) , im => to_ads_sfixed(0.889545)),
(re => to_ads_sfixed(-0.2724) , im => to_ads_sfixed(0.8816)),
(re => to_ads_sfixed(-0.27802) , im => to_ads_sfixed(0.873655)),
(re => to_ads_sfixed(-0.28364) , im => to_ads_sfixed(0.86571)),
(re => to_ads_sfixed(-0.28926) , im => to_ads_sfixed(0.857765)),
(re => to_ads_sfixed(-0.29488) , im => to_ads_sfixed(0.84982)),
(re => to_ads_sfixed(-0.3005) , im => to_ads_sfixed(0.841875)),
(re => to_ads_sfixed(-0.30612) , im => to_ads_sfixed(0.83393)),
(re => to_ads_sfixed(-0.31174) , im => to_ads_sfixed(0.825985)),
(re => to_ads_sfixed(-0.31736) , im => to_ads_sfixed(0.81804)),
(re => to_ads_sfixed(-0.32298) , im => to_ads_sfixed(0.810095)),
(re => to_ads_sfixed(-0.3286) , im => to_ads_sfixed(0.80215)),
(re => to_ads_sfixed(-0.33422) , im => to_ads_sfixed(0.794205)),
(re => to_ads_sfixed(-0.33984) , im => to_ads_sfixed(0.78626)),
(re => to_ads_sfixed(-0.34546) , im => to_ads_sfixed(0.778315)),
(re => to_ads_sfixed(-0.35108) , im => to_ads_sfixed(0.77037)),
(re => to_ads_sfixed(-0.3567) , im => to_ads_sfixed(0.762425)),
(re => to_ads_sfixed(-0.36232) , im => to_ads_sfixed(0.75448)),
(re => to_ads_sfixed(-0.36794) , im => to_ads_sfixed(0.746535)),
(re => to_ads_sfixed(-0.37356) , im => to_ads_sfixed(0.73859)),
(re => to_ads_sfixed(-0.37918) , im => to_ads_sfixed(0.730645)),
(re => to_ads_sfixed(-0.3848) , im => to_ads_sfixed(0.7227)),
(re => to_ads_sfixed(-0.39042) , im => to_ads_sfixed(0.714755)),
(re => to_ads_sfixed(-0.39604) , im => to_ads_sfixed(0.70681)),
(re => to_ads_sfixed(-0.40166) , im => to_ads_sfixed(0.698865)),
(re => to_ads_sfixed(-0.40728) , im => to_ads_sfixed(0.69092)),
(re => to_ads_sfixed(-0.4129) , im => to_ads_sfixed(0.682975)),
(re => to_ads_sfixed(-0.41852) , im => to_ads_sfixed(0.67503)),
(re => to_ads_sfixed(-0.42414) , im => to_ads_sfixed(0.667085)),
(re => to_ads_sfixed(-0.42976) , im => to_ads_sfixed(0.65914)),
(re => to_ads_sfixed(-0.43538) , im => to_ads_sfixed(0.651195)),
(re => to_ads_sfixed(-0.441) , im => to_ads_sfixed(0.64325)),
(re => to_ads_sfixed(-0.44662) , im => to_ads_sfixed(0.635305)),
(re => to_ads_sfixed(-0.45224) , im => to_ads_sfixed(0.62736)),
(re => to_ads_sfixed(-0.45786) , im => to_ads_sfixed(0.619415)),
(re => to_ads_sfixed(-0.46348) , im => to_ads_sfixed(0.61147)),
(re => to_ads_sfixed(-0.4691) , im => to_ads_sfixed(0.603525)),
(re => to_ads_sfixed(-0.47472) , im => to_ads_sfixed(0.59558)),
(re => to_ads_sfixed(-0.48034) , im => to_ads_sfixed(0.587635)),
(re => to_ads_sfixed(-0.48596) , im => to_ads_sfixed(0.57969)),
(re => to_ads_sfixed(-0.49158) , im => to_ads_sfixed(0.571745)),
(re => to_ads_sfixed(-0.4972) , im => to_ads_sfixed(0.5638)),
(re => to_ads_sfixed(-0.50282) , im => to_ads_sfixed(0.555855)),
(re => to_ads_sfixed(-0.50844) , im => to_ads_sfixed(0.54791)),
(re => to_ads_sfixed(-0.51406) , im => to_ads_sfixed(0.539965)),
(re => to_ads_sfixed(-0.51968) , im => to_ads_sfixed(0.53202)),
(re => to_ads_sfixed(-0.5253) , im => to_ads_sfixed(0.524075)),
(re => to_ads_sfixed(-0.53092) , im => to_ads_sfixed(0.51613)),
(re => to_ads_sfixed(-0.53654) , im => to_ads_sfixed(0.508185)),
(re => to_ads_sfixed(-0.54216) , im => to_ads_sfixed(0.50024)),
(re => to_ads_sfixed(-0.54778) , im => to_ads_sfixed(0.492295)),
(re => to_ads_sfixed(-0.5534) , im => to_ads_sfixed(0.48435)),
(re => to_ads_sfixed(-0.55902) , im => to_ads_sfixed(0.476405)),
(re => to_ads_sfixed(-0.56464) , im => to_ads_sfixed(0.46846)),
(re => to_ads_sfixed(-0.57026) , im => to_ads_sfixed(0.460515)),
(re => to_ads_sfixed(-0.57588) , im => to_ads_sfixed(0.45257)),
(re => to_ads_sfixed(-0.5815) , im => to_ads_sfixed(0.444625)),
(re => to_ads_sfixed(-0.58712) , im => to_ads_sfixed(0.43668)),
(re => to_ads_sfixed(-0.59274) , im => to_ads_sfixed(0.428735)),
(re => to_ads_sfixed(-0.59836) , im => to_ads_sfixed(0.42079)),
(re => to_ads_sfixed(-0.60398) , im => to_ads_sfixed(0.412845)),
(re => to_ads_sfixed(-0.6096) , im => to_ads_sfixed(0.4049)),
(re => to_ads_sfixed(-0.61522) , im => to_ads_sfixed(0.396955)),
(re => to_ads_sfixed(-0.62084) , im => to_ads_sfixed(0.38901)),
(re => to_ads_sfixed(-0.62646) , im => to_ads_sfixed(0.381065)),
(re => to_ads_sfixed(-0.63208) , im => to_ads_sfixed(0.37312)),
(re => to_ads_sfixed(-0.6377) , im => to_ads_sfixed(0.365175)),
(re => to_ads_sfixed(-0.64332) , im => to_ads_sfixed(0.35723)),
(re => to_ads_sfixed(-0.64894) , im => to_ads_sfixed(0.349285)),
(re => to_ads_sfixed(-0.65456) , im => to_ads_sfixed(0.34134)),
(re => to_ads_sfixed(-0.66018) , im => to_ads_sfixed(0.333395)),
(re => to_ads_sfixed(-0.6658) , im => to_ads_sfixed(0.32545)),
(re => to_ads_sfixed(-0.67142) , im => to_ads_sfixed(0.317505)),
(re => to_ads_sfixed(-0.67704) , im => to_ads_sfixed(0.30956)),
(re => to_ads_sfixed(-0.68266) , im => to_ads_sfixed(0.301615)),
(re => to_ads_sfixed(-0.68828) , im => to_ads_sfixed(0.29367)),
(re => to_ads_sfixed(-0.6939) , im => to_ads_sfixed(0.285725)),
(re => to_ads_sfixed(-0.69952) , im => to_ads_sfixed(0.27778)),
(re => to_ads_sfixed(-0.70514) , im => to_ads_sfixed(0.269835)),
(re => to_ads_sfixed(-0.71076) , im => to_ads_sfixed(0.26189)),
(re => to_ads_sfixed(-0.71638) , im => to_ads_sfixed(0.253945)),
(re => to_ads_sfixed(-0.722) , im => to_ads_sfixed(0.246)),
(re => to_ads_sfixed(-0.7222329) , im => to_ads_sfixed(0.24467075)),
(re => to_ads_sfixed(-0.7224658) , im => to_ads_sfixed(0.2433415)),
(re => to_ads_sfixed(-0.7226987) , im => to_ads_sfixed(0.24201225)),
(re => to_ads_sfixed(-0.7229316) , im => to_ads_sfixed(0.240683)),
(re => to_ads_sfixed(-0.7231645) , im => to_ads_sfixed(0.23935375)),
(re => to_ads_sfixed(-0.7233974) , im => to_ads_sfixed(0.2380245)),
(re => to_ads_sfixed(-0.7236303) , im => to_ads_sfixed(0.23669525)),
(re => to_ads_sfixed(-0.7238632) , im => to_ads_sfixed(0.235366)),
(re => to_ads_sfixed(-0.7240961) , im => to_ads_sfixed(0.23403675)),
(re => to_ads_sfixed(-0.724329) , im => to_ads_sfixed(0.2327075)),
(re => to_ads_sfixed(-0.7245619) , im => to_ads_sfixed(0.23137825)),
(re => to_ads_sfixed(-0.7247948) , im => to_ads_sfixed(0.230049)),
(re => to_ads_sfixed(-0.7250277) , im => to_ads_sfixed(0.22871975)),
(re => to_ads_sfixed(-0.7252606) , im => to_ads_sfixed(0.2273905)),
(re => to_ads_sfixed(-0.7254935) , im => to_ads_sfixed(0.22606125)),
(re => to_ads_sfixed(-0.7257264) , im => to_ads_sfixed(0.224732)),
(re => to_ads_sfixed(-0.7259593) , im => to_ads_sfixed(0.22340275)),
(re => to_ads_sfixed(-0.7261922) , im => to_ads_sfixed(0.2220735)),
(re => to_ads_sfixed(-0.7264251) , im => to_ads_sfixed(0.22074425)),
(re => to_ads_sfixed(-0.726658) , im => to_ads_sfixed(0.219415)),
(re => to_ads_sfixed(-0.7268909) , im => to_ads_sfixed(0.21808575)),
(re => to_ads_sfixed(-0.7271238) , im => to_ads_sfixed(0.2167565)),
(re => to_ads_sfixed(-0.7273567) , im => to_ads_sfixed(0.21542725)),
(re => to_ads_sfixed(-0.7275896) , im => to_ads_sfixed(0.214098)),
(re => to_ads_sfixed(-0.7278225) , im => to_ads_sfixed(0.21276875)),
(re => to_ads_sfixed(-0.7280554) , im => to_ads_sfixed(0.2114395)),
(re => to_ads_sfixed(-0.7282883) , im => to_ads_sfixed(0.21011025)),
(re => to_ads_sfixed(-0.7285212) , im => to_ads_sfixed(0.208781)),
(re => to_ads_sfixed(-0.7287541) , im => to_ads_sfixed(0.20745175)),
(re => to_ads_sfixed(-0.728987) , im => to_ads_sfixed(0.2061225)),
(re => to_ads_sfixed(-0.7292199) , im => to_ads_sfixed(0.20479325)),
(re => to_ads_sfixed(-0.7294528) , im => to_ads_sfixed(0.203464)),
(re => to_ads_sfixed(-0.7296857) , im => to_ads_sfixed(0.20213475)),
(re => to_ads_sfixed(-0.7299186) , im => to_ads_sfixed(0.2008055)),
(re => to_ads_sfixed(-0.7301515) , im => to_ads_sfixed(0.19947625)),
(re => to_ads_sfixed(-0.7303844) , im => to_ads_sfixed(0.198147)),
(re => to_ads_sfixed(-0.7306173) , im => to_ads_sfixed(0.19681775)),
(re => to_ads_sfixed(-0.7308502) , im => to_ads_sfixed(0.1954885)),
(re => to_ads_sfixed(-0.7310831) , im => to_ads_sfixed(0.19415925)),
(re => to_ads_sfixed(-0.731316) , im => to_ads_sfixed(0.19283)),
(re => to_ads_sfixed(-0.7315489) , im => to_ads_sfixed(0.19150075)),
(re => to_ads_sfixed(-0.7317818) , im => to_ads_sfixed(0.1901715)),
(re => to_ads_sfixed(-0.7320147) , im => to_ads_sfixed(0.18884225)),
(re => to_ads_sfixed(-0.7322476) , im => to_ads_sfixed(0.187513)),
(re => to_ads_sfixed(-0.7324805) , im => to_ads_sfixed(0.18618375)),
(re => to_ads_sfixed(-0.7327134) , im => to_ads_sfixed(0.1848545)),
(re => to_ads_sfixed(-0.7329463) , im => to_ads_sfixed(0.18352525)),
(re => to_ads_sfixed(-0.7331792) , im => to_ads_sfixed(0.182196)),
(re => to_ads_sfixed(-0.7334121) , im => to_ads_sfixed(0.18086675)),
(re => to_ads_sfixed(-0.733645) , im => to_ads_sfixed(0.1795375)),
(re => to_ads_sfixed(-0.7338779) , im => to_ads_sfixed(0.17820825)),
(re => to_ads_sfixed(-0.7341108) , im => to_ads_sfixed(0.176879)),
(re => to_ads_sfixed(-0.7343437) , im => to_ads_sfixed(0.17554975)),
(re => to_ads_sfixed(-0.7345766) , im => to_ads_sfixed(0.1742205)),
(re => to_ads_sfixed(-0.7348095) , im => to_ads_sfixed(0.17289125)),
(re => to_ads_sfixed(-0.7350424) , im => to_ads_sfixed(0.171562)),
(re => to_ads_sfixed(-0.7352753) , im => to_ads_sfixed(0.17023275)),
(re => to_ads_sfixed(-0.7355082) , im => to_ads_sfixed(0.1689035)),
(re => to_ads_sfixed(-0.7357411) , im => to_ads_sfixed(0.16757425)),
(re => to_ads_sfixed(-0.735974) , im => to_ads_sfixed(0.166245)),
(re => to_ads_sfixed(-0.7362069) , im => to_ads_sfixed(0.16491575)),
(re => to_ads_sfixed(-0.7364398) , im => to_ads_sfixed(0.1635865)),
(re => to_ads_sfixed(-0.7366727) , im => to_ads_sfixed(0.16225725)),
(re => to_ads_sfixed(-0.7369056) , im => to_ads_sfixed(0.160928)),
(re => to_ads_sfixed(-0.7371385) , im => to_ads_sfixed(0.15959875)),
(re => to_ads_sfixed(-0.7373714) , im => to_ads_sfixed(0.1582695)),
(re => to_ads_sfixed(-0.7376043) , im => to_ads_sfixed(0.15694025)),
(re => to_ads_sfixed(-0.7378372) , im => to_ads_sfixed(0.155611)),
(re => to_ads_sfixed(-0.7380701) , im => to_ads_sfixed(0.15428175)),
(re => to_ads_sfixed(-0.738303) , im => to_ads_sfixed(0.1529525)),
(re => to_ads_sfixed(-0.7385359) , im => to_ads_sfixed(0.15162325)),
(re => to_ads_sfixed(-0.7387688) , im => to_ads_sfixed(0.150294)),
(re => to_ads_sfixed(-0.7390017) , im => to_ads_sfixed(0.14896475)),
(re => to_ads_sfixed(-0.7392346) , im => to_ads_sfixed(0.1476355)),
(re => to_ads_sfixed(-0.7394675) , im => to_ads_sfixed(0.14630625)),
(re => to_ads_sfixed(-0.7397004) , im => to_ads_sfixed(0.144977)),
(re => to_ads_sfixed(-0.7399333) , im => to_ads_sfixed(0.14364775)),
(re => to_ads_sfixed(-0.7401662) , im => to_ads_sfixed(0.1423185)),
(re => to_ads_sfixed(-0.7403991) , im => to_ads_sfixed(0.14098925)),
(re => to_ads_sfixed(-0.740632) , im => to_ads_sfixed(0.13966)),
(re => to_ads_sfixed(-0.7408649) , im => to_ads_sfixed(0.13833075)),
(re => to_ads_sfixed(-0.7410978) , im => to_ads_sfixed(0.1370015)),
(re => to_ads_sfixed(-0.7413307) , im => to_ads_sfixed(0.13567225)),
(re => to_ads_sfixed(-0.7415636) , im => to_ads_sfixed(0.134343)),
(re => to_ads_sfixed(-0.7417965) , im => to_ads_sfixed(0.13301375)),
(re => to_ads_sfixed(-0.7420294) , im => to_ads_sfixed(0.1316845)),
(re => to_ads_sfixed(-0.7422623) , im => to_ads_sfixed(0.13035525)),
(re => to_ads_sfixed(-0.7424952) , im => to_ads_sfixed(0.129026)),
(re => to_ads_sfixed(-0.7427281) , im => to_ads_sfixed(0.12769675)),
(re => to_ads_sfixed(-0.742961) , im => to_ads_sfixed(0.1263675)),
(re => to_ads_sfixed(-0.7431939) , im => to_ads_sfixed(0.12503825)),
(re => to_ads_sfixed(-0.7434268) , im => to_ads_sfixed(0.123709)),
(re => to_ads_sfixed(-0.7436597) , im => to_ads_sfixed(0.12237975)),
(re => to_ads_sfixed(-0.7438926) , im => to_ads_sfixed(0.1210505)),
(re => to_ads_sfixed(-0.7441255) , im => to_ads_sfixed(0.11972125)),
(re => to_ads_sfixed(-0.7443584) , im => to_ads_sfixed(0.118392)),
(re => to_ads_sfixed(-0.7445913) , im => to_ads_sfixed(0.11706275)),
(re => to_ads_sfixed(-0.7448242) , im => to_ads_sfixed(0.1157335)),
(re => to_ads_sfixed(-0.7450571) , im => to_ads_sfixed(0.11440425)),
(re => to_ads_sfixed(-0.74529) , im => to_ads_sfixed(0.113075)),
(re => to_ads_sfixed(-0.7418371) , im => to_ads_sfixed(0.10604425)),
(re => to_ads_sfixed(-0.7383842) , im => to_ads_sfixed(0.0990135)),
(re => to_ads_sfixed(-0.7349313) , im => to_ads_sfixed(0.09198275)),
(re => to_ads_sfixed(-0.7314784) , im => to_ads_sfixed(0.084952)),
(re => to_ads_sfixed(-0.7280255) , im => to_ads_sfixed(0.07792125)),
(re => to_ads_sfixed(-0.7245726) , im => to_ads_sfixed(0.0708905)),
(re => to_ads_sfixed(-0.7211197) , im => to_ads_sfixed(0.06385975)),
(re => to_ads_sfixed(-0.7176668) , im => to_ads_sfixed(0.056829)),
(re => to_ads_sfixed(-0.7142139) , im => to_ads_sfixed(0.04979825)),
(re => to_ads_sfixed(-0.710761) , im => to_ads_sfixed(0.0427675)),
(re => to_ads_sfixed(-0.7073081) , im => to_ads_sfixed(0.03573675)),
(re => to_ads_sfixed(-0.7038552) , im => to_ads_sfixed(0.028706)),
(re => to_ads_sfixed(-0.7004023) , im => to_ads_sfixed(0.02167525)),
(re => to_ads_sfixed(-0.6969494) , im => to_ads_sfixed(0.0146445)),
(re => to_ads_sfixed(-0.6934965) , im => to_ads_sfixed(0.00761375)),
(re => to_ads_sfixed(-0.6900436) , im => to_ads_sfixed(0.000583)),
(re => to_ads_sfixed(-0.6865907) , im => to_ads_sfixed(-0.00644775)),
(re => to_ads_sfixed(-0.6831378) , im => to_ads_sfixed(-0.0134785)),
(re => to_ads_sfixed(-0.6796849) , im => to_ads_sfixed(-0.02050925)),
(re => to_ads_sfixed(-0.676232) , im => to_ads_sfixed(-0.02754)),
(re => to_ads_sfixed(-0.6727791) , im => to_ads_sfixed(-0.03457075)),
(re => to_ads_sfixed(-0.6693262) , im => to_ads_sfixed(-0.0416015)),
(re => to_ads_sfixed(-0.6658733) , im => to_ads_sfixed(-0.04863225)),
(re => to_ads_sfixed(-0.6624204) , im => to_ads_sfixed(-0.055663)),
(re => to_ads_sfixed(-0.6589675) , im => to_ads_sfixed(-0.06269375)),
(re => to_ads_sfixed(-0.6555146) , im => to_ads_sfixed(-0.0697245)),
(re => to_ads_sfixed(-0.6520617) , im => to_ads_sfixed(-0.07675525)),
(re => to_ads_sfixed(-0.6486088) , im => to_ads_sfixed(-0.083786)),
(re => to_ads_sfixed(-0.6451559) , im => to_ads_sfixed(-0.09081675)),
(re => to_ads_sfixed(-0.641703) , im => to_ads_sfixed(-0.0978475)),
(re => to_ads_sfixed(-0.6382501) , im => to_ads_sfixed(-0.10487825)),
(re => to_ads_sfixed(-0.6347972) , im => to_ads_sfixed(-0.111909)),
(re => to_ads_sfixed(-0.6313443) , im => to_ads_sfixed(-0.11893975)),
(re => to_ads_sfixed(-0.6278914) , im => to_ads_sfixed(-0.1259705)),
(re => to_ads_sfixed(-0.6244385) , im => to_ads_sfixed(-0.13300125)),
(re => to_ads_sfixed(-0.6209856) , im => to_ads_sfixed(-0.140032)),
(re => to_ads_sfixed(-0.6175327) , im => to_ads_sfixed(-0.14706275)),
(re => to_ads_sfixed(-0.6140798) , im => to_ads_sfixed(-0.1540935)),
(re => to_ads_sfixed(-0.6106269) , im => to_ads_sfixed(-0.16112425)),
(re => to_ads_sfixed(-0.607174) , im => to_ads_sfixed(-0.168155)),
(re => to_ads_sfixed(-0.6037211) , im => to_ads_sfixed(-0.17518575)),
(re => to_ads_sfixed(-0.6002682) , im => to_ads_sfixed(-0.1822165)),
(re => to_ads_sfixed(-0.5968153) , im => to_ads_sfixed(-0.18924725)),
(re => to_ads_sfixed(-0.5933624) , im => to_ads_sfixed(-0.196278)),
(re => to_ads_sfixed(-0.5899095) , im => to_ads_sfixed(-0.20330875)),
(re => to_ads_sfixed(-0.5864566) , im => to_ads_sfixed(-0.2103395)),
(re => to_ads_sfixed(-0.5830037) , im => to_ads_sfixed(-0.21737025)),
(re => to_ads_sfixed(-0.5795508) , im => to_ads_sfixed(-0.224401)),
(re => to_ads_sfixed(-0.5760979) , im => to_ads_sfixed(-0.23143175)),
(re => to_ads_sfixed(-0.572645) , im => to_ads_sfixed(-0.2384625)),
(re => to_ads_sfixed(-0.5691921) , im => to_ads_sfixed(-0.24549325)),
(re => to_ads_sfixed(-0.5657392) , im => to_ads_sfixed(-0.252524)),
(re => to_ads_sfixed(-0.5622863) , im => to_ads_sfixed(-0.25955475)),
(re => to_ads_sfixed(-0.5588334) , im => to_ads_sfixed(-0.2665855)),
(re => to_ads_sfixed(-0.5553805) , im => to_ads_sfixed(-0.27361625)),
(re => to_ads_sfixed(-0.5519276) , im => to_ads_sfixed(-0.280647)),
(re => to_ads_sfixed(-0.5484747) , im => to_ads_sfixed(-0.28767775)),
(re => to_ads_sfixed(-0.5450218) , im => to_ads_sfixed(-0.2947085)),
(re => to_ads_sfixed(-0.5415689) , im => to_ads_sfixed(-0.30173925)),
(re => to_ads_sfixed(-0.538116) , im => to_ads_sfixed(-0.30877)),
(re => to_ads_sfixed(-0.5346631) , im => to_ads_sfixed(-0.31580075)),
(re => to_ads_sfixed(-0.5312102) , im => to_ads_sfixed(-0.3228315)),
(re => to_ads_sfixed(-0.5277573) , im => to_ads_sfixed(-0.32986225)),
(re => to_ads_sfixed(-0.5243044) , im => to_ads_sfixed(-0.336893)),
(re => to_ads_sfixed(-0.5208515) , im => to_ads_sfixed(-0.34392375)),
(re => to_ads_sfixed(-0.5173986) , im => to_ads_sfixed(-0.3509545)),
(re => to_ads_sfixed(-0.5139457) , im => to_ads_sfixed(-0.35798525)),
(re => to_ads_sfixed(-0.5104928) , im => to_ads_sfixed(-0.365016)),
(re => to_ads_sfixed(-0.5070399) , im => to_ads_sfixed(-0.37204675)),
(re => to_ads_sfixed(-0.503587) , im => to_ads_sfixed(-0.3790775)),
(re => to_ads_sfixed(-0.5001341) , im => to_ads_sfixed(-0.38610825)),
(re => to_ads_sfixed(-0.4966812) , im => to_ads_sfixed(-0.393139)),
(re => to_ads_sfixed(-0.4932283) , im => to_ads_sfixed(-0.40016975)),
(re => to_ads_sfixed(-0.4897754) , im => to_ads_sfixed(-0.4072005)),
(re => to_ads_sfixed(-0.4863225) , im => to_ads_sfixed(-0.41423125)),
(re => to_ads_sfixed(-0.4828696) , im => to_ads_sfixed(-0.421262)),
(re => to_ads_sfixed(-0.4794167) , im => to_ads_sfixed(-0.42829275)),
(re => to_ads_sfixed(-0.4759638) , im => to_ads_sfixed(-0.4353235)),
(re => to_ads_sfixed(-0.4725109) , im => to_ads_sfixed(-0.44235425)),
(re => to_ads_sfixed(-0.469058) , im => to_ads_sfixed(-0.449385)),
(re => to_ads_sfixed(-0.4656051) , im => to_ads_sfixed(-0.45641575)),
(re => to_ads_sfixed(-0.4621522) , im => to_ads_sfixed(-0.4634465)),
(re => to_ads_sfixed(-0.4586993) , im => to_ads_sfixed(-0.47047725)),
(re => to_ads_sfixed(-0.4552464) , im => to_ads_sfixed(-0.477508)),
(re => to_ads_sfixed(-0.4517935) , im => to_ads_sfixed(-0.48453875)),
(re => to_ads_sfixed(-0.4483406) , im => to_ads_sfixed(-0.4915695)),
(re => to_ads_sfixed(-0.4448877) , im => to_ads_sfixed(-0.49860025)),
(re => to_ads_sfixed(-0.4414348) , im => to_ads_sfixed(-0.505631)),
(re => to_ads_sfixed(-0.4379819) , im => to_ads_sfixed(-0.51266175)),
(re => to_ads_sfixed(-0.434529) , im => to_ads_sfixed(-0.5196925)),
(re => to_ads_sfixed(-0.4310761) , im => to_ads_sfixed(-0.52672325)),
(re => to_ads_sfixed(-0.4276232) , im => to_ads_sfixed(-0.533754)),
(re => to_ads_sfixed(-0.4241703) , im => to_ads_sfixed(-0.54078475)),
(re => to_ads_sfixed(-0.4207174) , im => to_ads_sfixed(-0.5478155)),
(re => to_ads_sfixed(-0.4172645) , im => to_ads_sfixed(-0.55484625)),
(re => to_ads_sfixed(-0.4138116) , im => to_ads_sfixed(-0.561877)),
(re => to_ads_sfixed(-0.4103587) , im => to_ads_sfixed(-0.56890775)),
(re => to_ads_sfixed(-0.4069058) , im => to_ads_sfixed(-0.5759385)),
(re => to_ads_sfixed(-0.4034529) , im => to_ads_sfixed(-0.58296925)),
(re => to_ads_sfixed(-0.4) , im => to_ads_sfixed(-0.59)),
(re => to_ads_sfixed(-0.39244466) , im => to_ads_sfixed(-0.58747292)),
(re => to_ads_sfixed(-0.38488932) , im => to_ads_sfixed(-0.58494584)),
(re => to_ads_sfixed(-0.37733398) , im => to_ads_sfixed(-0.58241876)),
(re => to_ads_sfixed(-0.36977864) , im => to_ads_sfixed(-0.57989168)),
(re => to_ads_sfixed(-0.3622233) , im => to_ads_sfixed(-0.5773646)),
(re => to_ads_sfixed(-0.35466796) , im => to_ads_sfixed(-0.57483752)),
(re => to_ads_sfixed(-0.34711262) , im => to_ads_sfixed(-0.57231044)),
(re => to_ads_sfixed(-0.33955728) , im => to_ads_sfixed(-0.56978336)),
(re => to_ads_sfixed(-0.33200194) , im => to_ads_sfixed(-0.56725628)),
(re => to_ads_sfixed(-0.3244466) , im => to_ads_sfixed(-0.5647292)),
(re => to_ads_sfixed(-0.31689126) , im => to_ads_sfixed(-0.56220212)),
(re => to_ads_sfixed(-0.30933592) , im => to_ads_sfixed(-0.55967504)),
(re => to_ads_sfixed(-0.30178058) , im => to_ads_sfixed(-0.55714796)),
(re => to_ads_sfixed(-0.29422524) , im => to_ads_sfixed(-0.55462088)),
(re => to_ads_sfixed(-0.2866699) , im => to_ads_sfixed(-0.5520938)),
(re => to_ads_sfixed(-0.27911456) , im => to_ads_sfixed(-0.54956672)),
(re => to_ads_sfixed(-0.27155922) , im => to_ads_sfixed(-0.54703964)),
(re => to_ads_sfixed(-0.26400388) , im => to_ads_sfixed(-0.54451256)),
(re => to_ads_sfixed(-0.25644854) , im => to_ads_sfixed(-0.54198548)),
(re => to_ads_sfixed(-0.2488932) , im => to_ads_sfixed(-0.5394584)),
(re => to_ads_sfixed(-0.24133786) , im => to_ads_sfixed(-0.53693132)),
(re => to_ads_sfixed(-0.23378252) , im => to_ads_sfixed(-0.53440424)),
(re => to_ads_sfixed(-0.22622718) , im => to_ads_sfixed(-0.53187716)),
(re => to_ads_sfixed(-0.21867184) , im => to_ads_sfixed(-0.52935008)),
(re => to_ads_sfixed(-0.2111165) , im => to_ads_sfixed(-0.526823)),
(re => to_ads_sfixed(-0.20356116) , im => to_ads_sfixed(-0.52429592)),
(re => to_ads_sfixed(-0.19600582) , im => to_ads_sfixed(-0.52176884)),
(re => to_ads_sfixed(-0.18845048) , im => to_ads_sfixed(-0.51924176)),
(re => to_ads_sfixed(-0.18089514) , im => to_ads_sfixed(-0.51671468)),
(re => to_ads_sfixed(-0.1733398) , im => to_ads_sfixed(-0.5141876)),
(re => to_ads_sfixed(-0.16578446) , im => to_ads_sfixed(-0.51166052)),
(re => to_ads_sfixed(-0.15822912) , im => to_ads_sfixed(-0.50913344)),
(re => to_ads_sfixed(-0.15067378) , im => to_ads_sfixed(-0.50660636)),
(re => to_ads_sfixed(-0.14311844) , im => to_ads_sfixed(-0.50407928)),
(re => to_ads_sfixed(-0.1355631) , im => to_ads_sfixed(-0.5015522)),
(re => to_ads_sfixed(-0.12800776) , im => to_ads_sfixed(-0.49902512)),
(re => to_ads_sfixed(-0.12045242) , im => to_ads_sfixed(-0.49649804)),
(re => to_ads_sfixed(-0.11289708) , im => to_ads_sfixed(-0.49397096)),
(re => to_ads_sfixed(-0.10534174) , im => to_ads_sfixed(-0.49144388)),
(re => to_ads_sfixed(-0.0977864) , im => to_ads_sfixed(-0.4889168)),
(re => to_ads_sfixed(-0.09023106) , im => to_ads_sfixed(-0.48638972)),
(re => to_ads_sfixed(-0.08267572) , im => to_ads_sfixed(-0.48386264)),
(re => to_ads_sfixed(-0.07512038) , im => to_ads_sfixed(-0.48133556)),
(re => to_ads_sfixed(-0.06756504) , im => to_ads_sfixed(-0.47880848)),
(re => to_ads_sfixed(-0.0600097) , im => to_ads_sfixed(-0.4762814)),
(re => to_ads_sfixed(-0.05245436) , im => to_ads_sfixed(-0.47375432)),
(re => to_ads_sfixed(-0.04489902) , im => to_ads_sfixed(-0.47122724)),
(re => to_ads_sfixed(-0.03734368) , im => to_ads_sfixed(-0.46870016)),
(re => to_ads_sfixed(-0.02978834) , im => to_ads_sfixed(-0.46617308)),
(re => to_ads_sfixed(-0.022233) , im => to_ads_sfixed(-0.463646)),
(re => to_ads_sfixed(-0.01467766) , im => to_ads_sfixed(-0.46111892)),
(re => to_ads_sfixed(-0.00712232) , im => to_ads_sfixed(-0.45859184)),
(re => to_ads_sfixed(0.00043302) , im => to_ads_sfixed(-0.45606476)),
(re => to_ads_sfixed(0.00798836) , im => to_ads_sfixed(-0.45353768)),
(re => to_ads_sfixed(0.0155437) , im => to_ads_sfixed(-0.4510106)),
(re => to_ads_sfixed(0.02309904) , im => to_ads_sfixed(-0.44848352)),
(re => to_ads_sfixed(0.03065438) , im => to_ads_sfixed(-0.44595644)),
(re => to_ads_sfixed(0.03820972) , im => to_ads_sfixed(-0.44342936)),
(re => to_ads_sfixed(0.04576506) , im => to_ads_sfixed(-0.44090228)),
(re => to_ads_sfixed(0.0533204) , im => to_ads_sfixed(-0.4383752)),
(re => to_ads_sfixed(0.06087574) , im => to_ads_sfixed(-0.43584812)),
(re => to_ads_sfixed(0.06843108) , im => to_ads_sfixed(-0.43332104)),
(re => to_ads_sfixed(0.07598642) , im => to_ads_sfixed(-0.43079396)),
(re => to_ads_sfixed(0.08354176) , im => to_ads_sfixed(-0.42826688)),
(re => to_ads_sfixed(0.0910971) , im => to_ads_sfixed(-0.4257398)),
(re => to_ads_sfixed(0.09865244) , im => to_ads_sfixed(-0.42321272)),
(re => to_ads_sfixed(0.10620778) , im => to_ads_sfixed(-0.42068564)),
(re => to_ads_sfixed(0.11376312) , im => to_ads_sfixed(-0.41815856)),
(re => to_ads_sfixed(0.12131846) , im => to_ads_sfixed(-0.41563148)),
(re => to_ads_sfixed(0.1288738) , im => to_ads_sfixed(-0.4131044)),
(re => to_ads_sfixed(0.13642914) , im => to_ads_sfixed(-0.41057732)),
(re => to_ads_sfixed(0.14398448) , im => to_ads_sfixed(-0.40805024)),
(re => to_ads_sfixed(0.15153982) , im => to_ads_sfixed(-0.40552316)),
(re => to_ads_sfixed(0.15909516) , im => to_ads_sfixed(-0.40299608)),
(re => to_ads_sfixed(0.1666505) , im => to_ads_sfixed(-0.400469)),
(re => to_ads_sfixed(0.17420584) , im => to_ads_sfixed(-0.39794192)),
(re => to_ads_sfixed(0.18176118) , im => to_ads_sfixed(-0.39541484)),
(re => to_ads_sfixed(0.18931652) , im => to_ads_sfixed(-0.39288776)),
(re => to_ads_sfixed(0.19687186) , im => to_ads_sfixed(-0.39036068)),
(re => to_ads_sfixed(0.2044272) , im => to_ads_sfixed(-0.3878336)),
(re => to_ads_sfixed(0.21198254) , im => to_ads_sfixed(-0.38530652)),
(re => to_ads_sfixed(0.21953788) , im => to_ads_sfixed(-0.38277944)),
(re => to_ads_sfixed(0.22709322) , im => to_ads_sfixed(-0.38025236)),
(re => to_ads_sfixed(0.23464856) , im => to_ads_sfixed(-0.37772528)),
(re => to_ads_sfixed(0.2422039) , im => to_ads_sfixed(-0.3751982)),
(re => to_ads_sfixed(0.24975924) , im => to_ads_sfixed(-0.37267112)),
(re => to_ads_sfixed(0.25731458) , im => to_ads_sfixed(-0.37014404)),
(re => to_ads_sfixed(0.26486992) , im => to_ads_sfixed(-0.36761696)),
(re => to_ads_sfixed(0.27242526) , im => to_ads_sfixed(-0.36508988)),
(re => to_ads_sfixed(0.2799806) , im => to_ads_sfixed(-0.3625628)),
(re => to_ads_sfixed(0.28753594) , im => to_ads_sfixed(-0.36003572)),
(re => to_ads_sfixed(0.29509128) , im => to_ads_sfixed(-0.35750864)),
(re => to_ads_sfixed(0.30264662) , im => to_ads_sfixed(-0.35498156)),
(re => to_ads_sfixed(0.31020196) , im => to_ads_sfixed(-0.35245448)),
(re => to_ads_sfixed(0.3177573) , im => to_ads_sfixed(-0.3499274)),
(re => to_ads_sfixed(0.32531264) , im => to_ads_sfixed(-0.34740032)),
(re => to_ads_sfixed(0.33286798) , im => to_ads_sfixed(-0.34487324)),
(re => to_ads_sfixed(0.34042332) , im => to_ads_sfixed(-0.34234616)),
(re => to_ads_sfixed(0.34797866) , im => to_ads_sfixed(-0.33981908)),
(re => to_ads_sfixed(0.355534) , im => to_ads_sfixed(-0.337292)),
(re => to_ads_sfixed(0.35537866) , im => to_ads_sfixed(-0.33441908)),
(re => to_ads_sfixed(0.35522332) , im => to_ads_sfixed(-0.33154616)),
(re => to_ads_sfixed(0.35506798) , im => to_ads_sfixed(-0.32867324)),
(re => to_ads_sfixed(0.35491264) , im => to_ads_sfixed(-0.32580032)),
(re => to_ads_sfixed(0.3547573) , im => to_ads_sfixed(-0.3229274)),
(re => to_ads_sfixed(0.35460196) , im => to_ads_sfixed(-0.32005448)),
(re => to_ads_sfixed(0.35444662) , im => to_ads_sfixed(-0.31718156)),
(re => to_ads_sfixed(0.35429128) , im => to_ads_sfixed(-0.31430864)),
(re => to_ads_sfixed(0.35413594) , im => to_ads_sfixed(-0.31143572)),
(re => to_ads_sfixed(0.3539806) , im => to_ads_sfixed(-0.3085628)),
(re => to_ads_sfixed(0.35382526) , im => to_ads_sfixed(-0.30568988)),
(re => to_ads_sfixed(0.35366992) , im => to_ads_sfixed(-0.30281696)),
(re => to_ads_sfixed(0.35351458) , im => to_ads_sfixed(-0.29994404)),
(re => to_ads_sfixed(0.35335924) , im => to_ads_sfixed(-0.29707112)),
(re => to_ads_sfixed(0.3532039) , im => to_ads_sfixed(-0.2941982)),
(re => to_ads_sfixed(0.35304856) , im => to_ads_sfixed(-0.29132528)),
(re => to_ads_sfixed(0.35289322) , im => to_ads_sfixed(-0.28845236)),
(re => to_ads_sfixed(0.35273788) , im => to_ads_sfixed(-0.28557944)),
(re => to_ads_sfixed(0.35258254) , im => to_ads_sfixed(-0.28270652)),
(re => to_ads_sfixed(0.3524272) , im => to_ads_sfixed(-0.2798336)),
(re => to_ads_sfixed(0.35227186) , im => to_ads_sfixed(-0.27696068)),
(re => to_ads_sfixed(0.35211652) , im => to_ads_sfixed(-0.27408776)),
(re => to_ads_sfixed(0.35196118) , im => to_ads_sfixed(-0.27121484)),
(re => to_ads_sfixed(0.35180584) , im => to_ads_sfixed(-0.26834192)),
(re => to_ads_sfixed(0.3516505) , im => to_ads_sfixed(-0.265469)),
(re => to_ads_sfixed(0.35149516) , im => to_ads_sfixed(-0.26259608)),
(re => to_ads_sfixed(0.35133982) , im => to_ads_sfixed(-0.25972316)),
(re => to_ads_sfixed(0.35118448) , im => to_ads_sfixed(-0.25685024)),
(re => to_ads_sfixed(0.35102914) , im => to_ads_sfixed(-0.25397732)),
(re => to_ads_sfixed(0.3508738) , im => to_ads_sfixed(-0.2511044)),
(re => to_ads_sfixed(0.35071846) , im => to_ads_sfixed(-0.24823148)),
(re => to_ads_sfixed(0.35056312) , im => to_ads_sfixed(-0.24535856)),
(re => to_ads_sfixed(0.35040778) , im => to_ads_sfixed(-0.24248564)),
(re => to_ads_sfixed(0.35025244) , im => to_ads_sfixed(-0.23961272)),
(re => to_ads_sfixed(0.3500971) , im => to_ads_sfixed(-0.2367398)),
(re => to_ads_sfixed(0.34994176) , im => to_ads_sfixed(-0.23386688)),
(re => to_ads_sfixed(0.34978642) , im => to_ads_sfixed(-0.23099396)),
(re => to_ads_sfixed(0.34963108) , im => to_ads_sfixed(-0.22812104)),
(re => to_ads_sfixed(0.34947574) , im => to_ads_sfixed(-0.22524812)),
(re => to_ads_sfixed(0.3493204) , im => to_ads_sfixed(-0.2223752)),
(re => to_ads_sfixed(0.34916506) , im => to_ads_sfixed(-0.21950228)),
(re => to_ads_sfixed(0.34900972) , im => to_ads_sfixed(-0.21662936)),
(re => to_ads_sfixed(0.34885438) , im => to_ads_sfixed(-0.21375644)),
(re => to_ads_sfixed(0.34869904) , im => to_ads_sfixed(-0.21088352)),
(re => to_ads_sfixed(0.3485437) , im => to_ads_sfixed(-0.2080106)),
(re => to_ads_sfixed(0.34838836) , im => to_ads_sfixed(-0.20513768)),
(re => to_ads_sfixed(0.34823302) , im => to_ads_sfixed(-0.20226476)),
(re => to_ads_sfixed(0.34807768) , im => to_ads_sfixed(-0.19939184)),
(re => to_ads_sfixed(0.34792234) , im => to_ads_sfixed(-0.19651892)),
(re => to_ads_sfixed(0.347767) , im => to_ads_sfixed(-0.193646)),
(re => to_ads_sfixed(0.34761166) , im => to_ads_sfixed(-0.19077308)),
(re => to_ads_sfixed(0.34745632) , im => to_ads_sfixed(-0.18790016)),
(re => to_ads_sfixed(0.34730098) , im => to_ads_sfixed(-0.18502724)),
(re => to_ads_sfixed(0.34714564) , im => to_ads_sfixed(-0.18215432)),
(re => to_ads_sfixed(0.3469903) , im => to_ads_sfixed(-0.1792814)),
(re => to_ads_sfixed(0.34683496) , im => to_ads_sfixed(-0.17640848)),
(re => to_ads_sfixed(0.34667962) , im => to_ads_sfixed(-0.17353556)),
(re => to_ads_sfixed(0.34652428) , im => to_ads_sfixed(-0.17066264)),
(re => to_ads_sfixed(0.34636894) , im => to_ads_sfixed(-0.16778972)),
(re => to_ads_sfixed(0.3462136) , im => to_ads_sfixed(-0.1649168)),
(re => to_ads_sfixed(0.34605826) , im => to_ads_sfixed(-0.16204388)),
(re => to_ads_sfixed(0.34590292) , im => to_ads_sfixed(-0.15917096)),
(re => to_ads_sfixed(0.34574758) , im => to_ads_sfixed(-0.15629804)),
(re => to_ads_sfixed(0.34559224) , im => to_ads_sfixed(-0.15342512)),
(re => to_ads_sfixed(0.3454369) , im => to_ads_sfixed(-0.1505522)),
(re => to_ads_sfixed(0.34528156) , im => to_ads_sfixed(-0.14767928)),
(re => to_ads_sfixed(0.34512622) , im => to_ads_sfixed(-0.14480636)),
(re => to_ads_sfixed(0.34497088) , im => to_ads_sfixed(-0.14193344)),
(re => to_ads_sfixed(0.34481554) , im => to_ads_sfixed(-0.13906052)),
(re => to_ads_sfixed(0.3446602) , im => to_ads_sfixed(-0.1361876)),
(re => to_ads_sfixed(0.34450486) , im => to_ads_sfixed(-0.13331468)),
(re => to_ads_sfixed(0.34434952) , im => to_ads_sfixed(-0.13044176)),
(re => to_ads_sfixed(0.34419418) , im => to_ads_sfixed(-0.12756884)),
(re => to_ads_sfixed(0.34403884) , im => to_ads_sfixed(-0.12469592)),
(re => to_ads_sfixed(0.3438835) , im => to_ads_sfixed(-0.121823)),
(re => to_ads_sfixed(0.34372816) , im => to_ads_sfixed(-0.11895008)),
(re => to_ads_sfixed(0.34357282) , im => to_ads_sfixed(-0.11607716)),
(re => to_ads_sfixed(0.34341748) , im => to_ads_sfixed(-0.11320424)),
(re => to_ads_sfixed(0.34326214) , im => to_ads_sfixed(-0.11033132)),
(re => to_ads_sfixed(0.3431068) , im => to_ads_sfixed(-0.1074584)),
(re => to_ads_sfixed(0.34295146) , im => to_ads_sfixed(-0.10458548)),
(re => to_ads_sfixed(0.34279612) , im => to_ads_sfixed(-0.10171256)),
(re => to_ads_sfixed(0.34264078) , im => to_ads_sfixed(-0.09883964)),
(re => to_ads_sfixed(0.34248544) , im => to_ads_sfixed(-0.09596672)),
(re => to_ads_sfixed(0.3423301) , im => to_ads_sfixed(-0.0930938)),
(re => to_ads_sfixed(0.34217476) , im => to_ads_sfixed(-0.09022088)),
(re => to_ads_sfixed(0.34201942) , im => to_ads_sfixed(-0.08734796)),
(re => to_ads_sfixed(0.34186408) , im => to_ads_sfixed(-0.08447504)),
(re => to_ads_sfixed(0.34170874) , im => to_ads_sfixed(-0.08160212)),
(re => to_ads_sfixed(0.3415534) , im => to_ads_sfixed(-0.0787292)),
(re => to_ads_sfixed(0.34139806) , im => to_ads_sfixed(-0.07585628)),
(re => to_ads_sfixed(0.34124272) , im => to_ads_sfixed(-0.07298336)),
(re => to_ads_sfixed(0.34108738) , im => to_ads_sfixed(-0.07011044)),
(re => to_ads_sfixed(0.34093204) , im => to_ads_sfixed(-0.06723752)),
(re => to_ads_sfixed(0.3407767) , im => to_ads_sfixed(-0.0643646)),
(re => to_ads_sfixed(0.34062136) , im => to_ads_sfixed(-0.06149168)),
(re => to_ads_sfixed(0.34046602) , im => to_ads_sfixed(-0.05861876)),
(re => to_ads_sfixed(0.34031068) , im => to_ads_sfixed(-0.05574584)),
(re => to_ads_sfixed(0.34015534) , im => to_ads_sfixed(-0.05287292)),
(re => to_ads_sfixed(0.34) , im => to_ads_sfixed(-0.05)),
(re => to_ads_sfixed(0.3403) , im => to_ads_sfixed(-0.0485)),
(re => to_ads_sfixed(0.3406) , im => to_ads_sfixed(-0.047)),
(re => to_ads_sfixed(0.3409) , im => to_ads_sfixed(-0.0455)),
(re => to_ads_sfixed(0.3412) , im => to_ads_sfixed(-0.044)),
(re => to_ads_sfixed(0.3415) , im => to_ads_sfixed(-0.0425)),
(re => to_ads_sfixed(0.3418) , im => to_ads_sfixed(-0.041)),
(re => to_ads_sfixed(0.3421) , im => to_ads_sfixed(-0.0395)),
(re => to_ads_sfixed(0.3424) , im => to_ads_sfixed(-0.038)),
(re => to_ads_sfixed(0.3427) , im => to_ads_sfixed(-0.0365)),
(re => to_ads_sfixed(0.343) , im => to_ads_sfixed(-0.035)),
(re => to_ads_sfixed(0.3433) , im => to_ads_sfixed(-0.0335)),
(re => to_ads_sfixed(0.3436) , im => to_ads_sfixed(-0.032)),
(re => to_ads_sfixed(0.3439) , im => to_ads_sfixed(-0.0305)),
(re => to_ads_sfixed(0.3442) , im => to_ads_sfixed(-0.029)),
(re => to_ads_sfixed(0.3445) , im => to_ads_sfixed(-0.0275)),
(re => to_ads_sfixed(0.3448) , im => to_ads_sfixed(-0.026)),
(re => to_ads_sfixed(0.3451) , im => to_ads_sfixed(-0.0245)),
(re => to_ads_sfixed(0.3454) , im => to_ads_sfixed(-0.023)),
(re => to_ads_sfixed(0.3457) , im => to_ads_sfixed(-0.0215)),
(re => to_ads_sfixed(0.346) , im => to_ads_sfixed(-0.02)),
(re => to_ads_sfixed(0.3463) , im => to_ads_sfixed(-0.0185)),
(re => to_ads_sfixed(0.3466) , im => to_ads_sfixed(-0.017)),
(re => to_ads_sfixed(0.3469) , im => to_ads_sfixed(-0.0155)),
(re => to_ads_sfixed(0.3472) , im => to_ads_sfixed(-0.014)),
(re => to_ads_sfixed(0.3475) , im => to_ads_sfixed(-0.0125)),
(re => to_ads_sfixed(0.3478) , im => to_ads_sfixed(-0.011)),
(re => to_ads_sfixed(0.3481) , im => to_ads_sfixed(-0.0095)),
(re => to_ads_sfixed(0.3484) , im => to_ads_sfixed(-0.008)),
(re => to_ads_sfixed(0.3487) , im => to_ads_sfixed(-0.0065)),
(re => to_ads_sfixed(0.349) , im => to_ads_sfixed(-0.005)),
(re => to_ads_sfixed(0.3493) , im => to_ads_sfixed(-0.0035)),
(re => to_ads_sfixed(0.3496) , im => to_ads_sfixed(-0.002)),
(re => to_ads_sfixed(0.3499) , im => to_ads_sfixed(-0.0005)),
(re => to_ads_sfixed(0.3502) , im => to_ads_sfixed(0.001)),
(re => to_ads_sfixed(0.3505) , im => to_ads_sfixed(0.0025)),
(re => to_ads_sfixed(0.3508) , im => to_ads_sfixed(0.004)),
(re => to_ads_sfixed(0.3511) , im => to_ads_sfixed(0.0055)),
(re => to_ads_sfixed(0.3514) , im => to_ads_sfixed(0.007)),
(re => to_ads_sfixed(0.3517) , im => to_ads_sfixed(0.0085)),
(re => to_ads_sfixed(0.352) , im => to_ads_sfixed(0.01)),
(re => to_ads_sfixed(0.3523) , im => to_ads_sfixed(0.0115)),
(re => to_ads_sfixed(0.3526) , im => to_ads_sfixed(0.013)),
(re => to_ads_sfixed(0.3529) , im => to_ads_sfixed(0.0145)),
(re => to_ads_sfixed(0.3532) , im => to_ads_sfixed(0.016)),
(re => to_ads_sfixed(0.3535) , im => to_ads_sfixed(0.0175)),
(re => to_ads_sfixed(0.3538) , im => to_ads_sfixed(0.019)),
(re => to_ads_sfixed(0.3541) , im => to_ads_sfixed(0.0205)),
(re => to_ads_sfixed(0.3544) , im => to_ads_sfixed(0.022)),
(re => to_ads_sfixed(0.3547) , im => to_ads_sfixed(0.0235)),
(re => to_ads_sfixed(0.355) , im => to_ads_sfixed(0.025)),
(re => to_ads_sfixed(0.3553) , im => to_ads_sfixed(0.0265)),
(re => to_ads_sfixed(0.3556) , im => to_ads_sfixed(0.028)),
(re => to_ads_sfixed(0.3559) , im => to_ads_sfixed(0.0295)),
(re => to_ads_sfixed(0.3562) , im => to_ads_sfixed(0.031)),
(re => to_ads_sfixed(0.3565) , im => to_ads_sfixed(0.0325)),
(re => to_ads_sfixed(0.3568) , im => to_ads_sfixed(0.034)),
(re => to_ads_sfixed(0.3571) , im => to_ads_sfixed(0.0355)),
(re => to_ads_sfixed(0.3574) , im => to_ads_sfixed(0.037)),
(re => to_ads_sfixed(0.3577) , im => to_ads_sfixed(0.0385)),
(re => to_ads_sfixed(0.358) , im => to_ads_sfixed(0.04)),
(re => to_ads_sfixed(0.3583) , im => to_ads_sfixed(0.0415)),
(re => to_ads_sfixed(0.3586) , im => to_ads_sfixed(0.043)),
(re => to_ads_sfixed(0.3589) , im => to_ads_sfixed(0.0445)),
(re => to_ads_sfixed(0.3592) , im => to_ads_sfixed(0.046)),
(re => to_ads_sfixed(0.3595) , im => to_ads_sfixed(0.0475)),
(re => to_ads_sfixed(0.3598) , im => to_ads_sfixed(0.049)),
(re => to_ads_sfixed(0.3601) , im => to_ads_sfixed(0.0505)),
(re => to_ads_sfixed(0.3604) , im => to_ads_sfixed(0.052)),
(re => to_ads_sfixed(0.3607) , im => to_ads_sfixed(0.0535)),
(re => to_ads_sfixed(0.361) , im => to_ads_sfixed(0.055)),
(re => to_ads_sfixed(0.3613) , im => to_ads_sfixed(0.0565)),
(re => to_ads_sfixed(0.3616) , im => to_ads_sfixed(0.058)),
(re => to_ads_sfixed(0.3619) , im => to_ads_sfixed(0.0595)),
(re => to_ads_sfixed(0.3622) , im => to_ads_sfixed(0.061)),
(re => to_ads_sfixed(0.3625) , im => to_ads_sfixed(0.0625)),
(re => to_ads_sfixed(0.3628) , im => to_ads_sfixed(0.064)),
(re => to_ads_sfixed(0.3631) , im => to_ads_sfixed(0.0655)),
(re => to_ads_sfixed(0.3634) , im => to_ads_sfixed(0.067)),
(re => to_ads_sfixed(0.3637) , im => to_ads_sfixed(0.0685)),
(re => to_ads_sfixed(0.364) , im => to_ads_sfixed(0.07)),
(re => to_ads_sfixed(0.3643) , im => to_ads_sfixed(0.0715)),
(re => to_ads_sfixed(0.3646) , im => to_ads_sfixed(0.073)),
(re => to_ads_sfixed(0.3649) , im => to_ads_sfixed(0.0745)),
(re => to_ads_sfixed(0.3652) , im => to_ads_sfixed(0.076)),
(re => to_ads_sfixed(0.3655) , im => to_ads_sfixed(0.0775)),
(re => to_ads_sfixed(0.3658) , im => to_ads_sfixed(0.079)),
(re => to_ads_sfixed(0.3661) , im => to_ads_sfixed(0.0805)),
(re => to_ads_sfixed(0.3664) , im => to_ads_sfixed(0.082)),
(re => to_ads_sfixed(0.3667) , im => to_ads_sfixed(0.0835)),
(re => to_ads_sfixed(0.367) , im => to_ads_sfixed(0.085)),
(re => to_ads_sfixed(0.3673) , im => to_ads_sfixed(0.0865)),
(re => to_ads_sfixed(0.3676) , im => to_ads_sfixed(0.088)),
(re => to_ads_sfixed(0.3679) , im => to_ads_sfixed(0.0895)),
(re => to_ads_sfixed(0.3682) , im => to_ads_sfixed(0.091)),
(re => to_ads_sfixed(0.3685) , im => to_ads_sfixed(0.0925)),
(re => to_ads_sfixed(0.3688) , im => to_ads_sfixed(0.094)),
(re => to_ads_sfixed(0.3691) , im => to_ads_sfixed(0.0955)),
(re => to_ads_sfixed(0.3694) , im => to_ads_sfixed(0.097)),
(re => to_ads_sfixed(0.3697) , im => to_ads_sfixed(0.0985)),
(re => to_ads_sfixed(0.37) , im => to_ads_sfixed(0.1)),
(re => to_ads_sfixed(0.36985) , im => to_ads_sfixed(0.10255)),
(re => to_ads_sfixed(0.3697) , im => to_ads_sfixed(0.1051)),
(re => to_ads_sfixed(0.36955) , im => to_ads_sfixed(0.10765)),
(re => to_ads_sfixed(0.3694) , im => to_ads_sfixed(0.1102)),
(re => to_ads_sfixed(0.36925) , im => to_ads_sfixed(0.11275)),
(re => to_ads_sfixed(0.3691) , im => to_ads_sfixed(0.1153)),
(re => to_ads_sfixed(0.36895) , im => to_ads_sfixed(0.11785)),
(re => to_ads_sfixed(0.3688) , im => to_ads_sfixed(0.1204)),
(re => to_ads_sfixed(0.36865) , im => to_ads_sfixed(0.12295)),
(re => to_ads_sfixed(0.3685) , im => to_ads_sfixed(0.1255)),
(re => to_ads_sfixed(0.36835) , im => to_ads_sfixed(0.12805)),
(re => to_ads_sfixed(0.3682) , im => to_ads_sfixed(0.1306)),
(re => to_ads_sfixed(0.36805) , im => to_ads_sfixed(0.13315)),
(re => to_ads_sfixed(0.3679) , im => to_ads_sfixed(0.1357)),
(re => to_ads_sfixed(0.36775) , im => to_ads_sfixed(0.13825)),
(re => to_ads_sfixed(0.3676) , im => to_ads_sfixed(0.1408)),
(re => to_ads_sfixed(0.36745) , im => to_ads_sfixed(0.14335)),
(re => to_ads_sfixed(0.3673) , im => to_ads_sfixed(0.1459)),
(re => to_ads_sfixed(0.36715) , im => to_ads_sfixed(0.14845)),
(re => to_ads_sfixed(0.367) , im => to_ads_sfixed(0.151)),
(re => to_ads_sfixed(0.36685) , im => to_ads_sfixed(0.15355)),
(re => to_ads_sfixed(0.3667) , im => to_ads_sfixed(0.1561)),
(re => to_ads_sfixed(0.36655) , im => to_ads_sfixed(0.15865)),
(re => to_ads_sfixed(0.3664) , im => to_ads_sfixed(0.1612)),
(re => to_ads_sfixed(0.36625) , im => to_ads_sfixed(0.16375)),
(re => to_ads_sfixed(0.3661) , im => to_ads_sfixed(0.1663)),
(re => to_ads_sfixed(0.36595) , im => to_ads_sfixed(0.16885)),
(re => to_ads_sfixed(0.3658) , im => to_ads_sfixed(0.1714)),
(re => to_ads_sfixed(0.36565) , im => to_ads_sfixed(0.17395)),
(re => to_ads_sfixed(0.3655) , im => to_ads_sfixed(0.1765)),
(re => to_ads_sfixed(0.36535) , im => to_ads_sfixed(0.17905)),
(re => to_ads_sfixed(0.3652) , im => to_ads_sfixed(0.1816)),
(re => to_ads_sfixed(0.36505) , im => to_ads_sfixed(0.18415)),
(re => to_ads_sfixed(0.3649) , im => to_ads_sfixed(0.1867)),
(re => to_ads_sfixed(0.36475) , im => to_ads_sfixed(0.18925)),
(re => to_ads_sfixed(0.3646) , im => to_ads_sfixed(0.1918)),
(re => to_ads_sfixed(0.36445) , im => to_ads_sfixed(0.19435)),
(re => to_ads_sfixed(0.3643) , im => to_ads_sfixed(0.1969)),
(re => to_ads_sfixed(0.36415) , im => to_ads_sfixed(0.19945)),
(re => to_ads_sfixed(0.364) , im => to_ads_sfixed(0.202)),
(re => to_ads_sfixed(0.36385) , im => to_ads_sfixed(0.20455)),
(re => to_ads_sfixed(0.3637) , im => to_ads_sfixed(0.2071)),
(re => to_ads_sfixed(0.36355) , im => to_ads_sfixed(0.20965)),
(re => to_ads_sfixed(0.3634) , im => to_ads_sfixed(0.2122)),
(re => to_ads_sfixed(0.36325) , im => to_ads_sfixed(0.21475)),
(re => to_ads_sfixed(0.3631) , im => to_ads_sfixed(0.2173)),
(re => to_ads_sfixed(0.36295) , im => to_ads_sfixed(0.21985)),
(re => to_ads_sfixed(0.3628) , im => to_ads_sfixed(0.2224)),
(re => to_ads_sfixed(0.36265) , im => to_ads_sfixed(0.22495)),
(re => to_ads_sfixed(0.3625) , im => to_ads_sfixed(0.2275)),
(re => to_ads_sfixed(0.36235) , im => to_ads_sfixed(0.23005)),
(re => to_ads_sfixed(0.3622) , im => to_ads_sfixed(0.2326)),
(re => to_ads_sfixed(0.36205) , im => to_ads_sfixed(0.23515)),
(re => to_ads_sfixed(0.3619) , im => to_ads_sfixed(0.2377)),
(re => to_ads_sfixed(0.36175) , im => to_ads_sfixed(0.24025)),
(re => to_ads_sfixed(0.3616) , im => to_ads_sfixed(0.2428)),
(re => to_ads_sfixed(0.36145) , im => to_ads_sfixed(0.24535)),
(re => to_ads_sfixed(0.3613) , im => to_ads_sfixed(0.2479)),
(re => to_ads_sfixed(0.36115) , im => to_ads_sfixed(0.25045)),
(re => to_ads_sfixed(0.361) , im => to_ads_sfixed(0.253)),
(re => to_ads_sfixed(0.36085) , im => to_ads_sfixed(0.25555)),
(re => to_ads_sfixed(0.3607) , im => to_ads_sfixed(0.2581)),
(re => to_ads_sfixed(0.36055) , im => to_ads_sfixed(0.26065)),
(re => to_ads_sfixed(0.3604) , im => to_ads_sfixed(0.2632)),
(re => to_ads_sfixed(0.36025) , im => to_ads_sfixed(0.26575)),
(re => to_ads_sfixed(0.3601) , im => to_ads_sfixed(0.2683)),
(re => to_ads_sfixed(0.35995) , im => to_ads_sfixed(0.27085)),
(re => to_ads_sfixed(0.3598) , im => to_ads_sfixed(0.2734)),
(re => to_ads_sfixed(0.35965) , im => to_ads_sfixed(0.27595)),
(re => to_ads_sfixed(0.3595) , im => to_ads_sfixed(0.2785)),
(re => to_ads_sfixed(0.35935) , im => to_ads_sfixed(0.28105)),
(re => to_ads_sfixed(0.3592) , im => to_ads_sfixed(0.2836)),
(re => to_ads_sfixed(0.35905) , im => to_ads_sfixed(0.28615)),
(re => to_ads_sfixed(0.3589) , im => to_ads_sfixed(0.2887)),
(re => to_ads_sfixed(0.35875) , im => to_ads_sfixed(0.29125)),
(re => to_ads_sfixed(0.3586) , im => to_ads_sfixed(0.2938)),
(re => to_ads_sfixed(0.35845) , im => to_ads_sfixed(0.29635)),
(re => to_ads_sfixed(0.3583) , im => to_ads_sfixed(0.2989)),
(re => to_ads_sfixed(0.35815) , im => to_ads_sfixed(0.30145)),
(re => to_ads_sfixed(0.358) , im => to_ads_sfixed(0.304)),
(re => to_ads_sfixed(0.35785) , im => to_ads_sfixed(0.30655)),
(re => to_ads_sfixed(0.3577) , im => to_ads_sfixed(0.3091)),
(re => to_ads_sfixed(0.35755) , im => to_ads_sfixed(0.31165)),
(re => to_ads_sfixed(0.3574) , im => to_ads_sfixed(0.3142)),
(re => to_ads_sfixed(0.35725) , im => to_ads_sfixed(0.31675)),
(re => to_ads_sfixed(0.3571) , im => to_ads_sfixed(0.3193)),
(re => to_ads_sfixed(0.35695) , im => to_ads_sfixed(0.32185)),
(re => to_ads_sfixed(0.3568) , im => to_ads_sfixed(0.3244)),
(re => to_ads_sfixed(0.35665) , im => to_ads_sfixed(0.32695)),
(re => to_ads_sfixed(0.3565) , im => to_ads_sfixed(0.3295)),
(re => to_ads_sfixed(0.35635) , im => to_ads_sfixed(0.33205)),
(re => to_ads_sfixed(0.3562) , im => to_ads_sfixed(0.3346)),
(re => to_ads_sfixed(0.35605) , im => to_ads_sfixed(0.33715)),
(re => to_ads_sfixed(0.3559) , im => to_ads_sfixed(0.3397)),
(re => to_ads_sfixed(0.35575) , im => to_ads_sfixed(0.34225)),
(re => to_ads_sfixed(0.3556) , im => to_ads_sfixed(0.3448)),
(re => to_ads_sfixed(0.35545) , im => to_ads_sfixed(0.34735)),
(re => to_ads_sfixed(0.3553) , im => to_ads_sfixed(0.3499)),
(re => to_ads_sfixed(0.35515) , im => to_ads_sfixed(0.35245)),
(re => to_ads_sfixed(0.355) , im => to_ads_sfixed(0.355)),
(re => to_ads_sfixed(0.35685) , im => to_ads_sfixed(0.35685)),
(re => to_ads_sfixed(0.3587) , im => to_ads_sfixed(0.3587)),
(re => to_ads_sfixed(0.36055) , im => to_ads_sfixed(0.36055)),
(re => to_ads_sfixed(0.3624) , im => to_ads_sfixed(0.3624)),
(re => to_ads_sfixed(0.36425) , im => to_ads_sfixed(0.36425)),
(re => to_ads_sfixed(0.3661) , im => to_ads_sfixed(0.3661)),
(re => to_ads_sfixed(0.36795) , im => to_ads_sfixed(0.36795)),
(re => to_ads_sfixed(0.3698) , im => to_ads_sfixed(0.3698)),
(re => to_ads_sfixed(0.37165) , im => to_ads_sfixed(0.37165)),
(re => to_ads_sfixed(0.3735) , im => to_ads_sfixed(0.3735)),
(re => to_ads_sfixed(0.37535) , im => to_ads_sfixed(0.37535)),
(re => to_ads_sfixed(0.3772) , im => to_ads_sfixed(0.3772)),
(re => to_ads_sfixed(0.37905) , im => to_ads_sfixed(0.37905)),
(re => to_ads_sfixed(0.3809) , im => to_ads_sfixed(0.3809)),
(re => to_ads_sfixed(0.38275) , im => to_ads_sfixed(0.38275)),
(re => to_ads_sfixed(0.3846) , im => to_ads_sfixed(0.3846)),
(re => to_ads_sfixed(0.38645) , im => to_ads_sfixed(0.38645)),
(re => to_ads_sfixed(0.3883) , im => to_ads_sfixed(0.3883)),
(re => to_ads_sfixed(0.39015) , im => to_ads_sfixed(0.39015)),
(re => to_ads_sfixed(0.392) , im => to_ads_sfixed(0.392)),
(re => to_ads_sfixed(0.39385) , im => to_ads_sfixed(0.39385)),
(re => to_ads_sfixed(0.3957) , im => to_ads_sfixed(0.3957)),
(re => to_ads_sfixed(0.39755) , im => to_ads_sfixed(0.39755)),
(re => to_ads_sfixed(0.3994) , im => to_ads_sfixed(0.3994)),
(re => to_ads_sfixed(0.40125) , im => to_ads_sfixed(0.40125)),
(re => to_ads_sfixed(0.4031) , im => to_ads_sfixed(0.4031)),
(re => to_ads_sfixed(0.40495) , im => to_ads_sfixed(0.40495)),
(re => to_ads_sfixed(0.4068) , im => to_ads_sfixed(0.4068)),
(re => to_ads_sfixed(0.40865) , im => to_ads_sfixed(0.40865)),
(re => to_ads_sfixed(0.4105) , im => to_ads_sfixed(0.4105)),
(re => to_ads_sfixed(0.41235) , im => to_ads_sfixed(0.41235)),
(re => to_ads_sfixed(0.4142) , im => to_ads_sfixed(0.4142)),
(re => to_ads_sfixed(0.41605) , im => to_ads_sfixed(0.41605)),
(re => to_ads_sfixed(0.4179) , im => to_ads_sfixed(0.4179)),
(re => to_ads_sfixed(0.41975) , im => to_ads_sfixed(0.41975)),
(re => to_ads_sfixed(0.4216) , im => to_ads_sfixed(0.4216)),
(re => to_ads_sfixed(0.42345) , im => to_ads_sfixed(0.42345)),
(re => to_ads_sfixed(0.4253) , im => to_ads_sfixed(0.4253)),
(re => to_ads_sfixed(0.42715) , im => to_ads_sfixed(0.42715)),
(re => to_ads_sfixed(0.429) , im => to_ads_sfixed(0.429)),
(re => to_ads_sfixed(0.43085) , im => to_ads_sfixed(0.43085)),
(re => to_ads_sfixed(0.4327) , im => to_ads_sfixed(0.4327)),
(re => to_ads_sfixed(0.43455) , im => to_ads_sfixed(0.43455)),
(re => to_ads_sfixed(0.4364) , im => to_ads_sfixed(0.4364)),
(re => to_ads_sfixed(0.43825) , im => to_ads_sfixed(0.43825)),
(re => to_ads_sfixed(0.4401) , im => to_ads_sfixed(0.4401)),
(re => to_ads_sfixed(0.44195) , im => to_ads_sfixed(0.44195)),
(re => to_ads_sfixed(0.4438) , im => to_ads_sfixed(0.4438)),
(re => to_ads_sfixed(0.44565) , im => to_ads_sfixed(0.44565)),
(re => to_ads_sfixed(0.4475) , im => to_ads_sfixed(0.4475)),
(re => to_ads_sfixed(0.44935) , im => to_ads_sfixed(0.44935)),
(re => to_ads_sfixed(0.4512) , im => to_ads_sfixed(0.4512)),
(re => to_ads_sfixed(0.45305) , im => to_ads_sfixed(0.45305)),
(re => to_ads_sfixed(0.4549) , im => to_ads_sfixed(0.4549)),
(re => to_ads_sfixed(0.45675) , im => to_ads_sfixed(0.45675)),
(re => to_ads_sfixed(0.4586) , im => to_ads_sfixed(0.4586)),
(re => to_ads_sfixed(0.46045) , im => to_ads_sfixed(0.46045)),
(re => to_ads_sfixed(0.4623) , im => to_ads_sfixed(0.4623)),
(re => to_ads_sfixed(0.46415) , im => to_ads_sfixed(0.46415)),
(re => to_ads_sfixed(0.466) , im => to_ads_sfixed(0.466)),
(re => to_ads_sfixed(0.46785) , im => to_ads_sfixed(0.46785)),
(re => to_ads_sfixed(0.4697) , im => to_ads_sfixed(0.4697)),
(re => to_ads_sfixed(0.47155) , im => to_ads_sfixed(0.47155)),
(re => to_ads_sfixed(0.4734) , im => to_ads_sfixed(0.4734)),
(re => to_ads_sfixed(0.47525) , im => to_ads_sfixed(0.47525)),
(re => to_ads_sfixed(0.4771) , im => to_ads_sfixed(0.4771)),
(re => to_ads_sfixed(0.47895) , im => to_ads_sfixed(0.47895)),
(re => to_ads_sfixed(0.4808) , im => to_ads_sfixed(0.4808)),
(re => to_ads_sfixed(0.48265) , im => to_ads_sfixed(0.48265)),
(re => to_ads_sfixed(0.4845) , im => to_ads_sfixed(0.4845)),
(re => to_ads_sfixed(0.48635) , im => to_ads_sfixed(0.48635)),
(re => to_ads_sfixed(0.4882) , im => to_ads_sfixed(0.4882)),
(re => to_ads_sfixed(0.49005) , im => to_ads_sfixed(0.49005)),
(re => to_ads_sfixed(0.4919) , im => to_ads_sfixed(0.4919)),
(re => to_ads_sfixed(0.49375) , im => to_ads_sfixed(0.49375)),
(re => to_ads_sfixed(0.4956) , im => to_ads_sfixed(0.4956)),
(re => to_ads_sfixed(0.49745) , im => to_ads_sfixed(0.49745)),
(re => to_ads_sfixed(0.4993) , im => to_ads_sfixed(0.4993)),
(re => to_ads_sfixed(0.50115) , im => to_ads_sfixed(0.50115)),
(re => to_ads_sfixed(0.503) , im => to_ads_sfixed(0.503)),
(re => to_ads_sfixed(0.50485) , im => to_ads_sfixed(0.50485)),
(re => to_ads_sfixed(0.5067) , im => to_ads_sfixed(0.5067)),
(re => to_ads_sfixed(0.50855) , im => to_ads_sfixed(0.50855)),
(re => to_ads_sfixed(0.5104) , im => to_ads_sfixed(0.5104)),
(re => to_ads_sfixed(0.51225) , im => to_ads_sfixed(0.51225)),
(re => to_ads_sfixed(0.5141) , im => to_ads_sfixed(0.5141)),
(re => to_ads_sfixed(0.51595) , im => to_ads_sfixed(0.51595)),
(re => to_ads_sfixed(0.5178) , im => to_ads_sfixed(0.5178)),
(re => to_ads_sfixed(0.51965) , im => to_ads_sfixed(0.51965)),
(re => to_ads_sfixed(0.5215) , im => to_ads_sfixed(0.5215)),
(re => to_ads_sfixed(0.52335) , im => to_ads_sfixed(0.52335)),
(re => to_ads_sfixed(0.5252) , im => to_ads_sfixed(0.5252)),
(re => to_ads_sfixed(0.52705) , im => to_ads_sfixed(0.52705)),
(re => to_ads_sfixed(0.5289) , im => to_ads_sfixed(0.5289)),
(re => to_ads_sfixed(0.53075) , im => to_ads_sfixed(0.53075)),
(re => to_ads_sfixed(0.5326) , im => to_ads_sfixed(0.5326)),
(re => to_ads_sfixed(0.53445) , im => to_ads_sfixed(0.53445)),
(re => to_ads_sfixed(0.5363) , im => to_ads_sfixed(0.5363)),
(re => to_ads_sfixed(0.53815) , im => to_ads_sfixed(0.53815)),
(re => to_ads_sfixed(0.54) , im => to_ads_sfixed(0.54)),
(re => to_ads_sfixed(0.5346) , im => to_ads_sfixed(0.5426)),
(re => to_ads_sfixed(0.5292) , im => to_ads_sfixed(0.5452)),
(re => to_ads_sfixed(0.5238) , im => to_ads_sfixed(0.5478)),
(re => to_ads_sfixed(0.5184) , im => to_ads_sfixed(0.5504)),
(re => to_ads_sfixed(0.513) , im => to_ads_sfixed(0.553)),
(re => to_ads_sfixed(0.5076) , im => to_ads_sfixed(0.5556)),
(re => to_ads_sfixed(0.5022) , im => to_ads_sfixed(0.5582)),
(re => to_ads_sfixed(0.4968) , im => to_ads_sfixed(0.5608)),
(re => to_ads_sfixed(0.4914) , im => to_ads_sfixed(0.5634)),
(re => to_ads_sfixed(0.486) , im => to_ads_sfixed(0.566)),
(re => to_ads_sfixed(0.4806) , im => to_ads_sfixed(0.5686)),
(re => to_ads_sfixed(0.4752) , im => to_ads_sfixed(0.5712)),
(re => to_ads_sfixed(0.4698) , im => to_ads_sfixed(0.5738)),
(re => to_ads_sfixed(0.4644) , im => to_ads_sfixed(0.5764)),
(re => to_ads_sfixed(0.459) , im => to_ads_sfixed(0.579)),
(re => to_ads_sfixed(0.4536) , im => to_ads_sfixed(0.5816)),
(re => to_ads_sfixed(0.4482) , im => to_ads_sfixed(0.5842)),
(re => to_ads_sfixed(0.4428) , im => to_ads_sfixed(0.5868)),
(re => to_ads_sfixed(0.4374) , im => to_ads_sfixed(0.5894)),
(re => to_ads_sfixed(0.432) , im => to_ads_sfixed(0.592)),
(re => to_ads_sfixed(0.4266) , im => to_ads_sfixed(0.5946)),
(re => to_ads_sfixed(0.4212) , im => to_ads_sfixed(0.5972)),
(re => to_ads_sfixed(0.4158) , im => to_ads_sfixed(0.5998)),
(re => to_ads_sfixed(0.4104) , im => to_ads_sfixed(0.6024)),
(re => to_ads_sfixed(0.405) , im => to_ads_sfixed(0.605)),
(re => to_ads_sfixed(0.3996) , im => to_ads_sfixed(0.6076)),
(re => to_ads_sfixed(0.3942) , im => to_ads_sfixed(0.6102)),
(re => to_ads_sfixed(0.3888) , im => to_ads_sfixed(0.6128)),
(re => to_ads_sfixed(0.3834) , im => to_ads_sfixed(0.6154)),
(re => to_ads_sfixed(0.378) , im => to_ads_sfixed(0.618)),
(re => to_ads_sfixed(0.3726) , im => to_ads_sfixed(0.6206)),
(re => to_ads_sfixed(0.3672) , im => to_ads_sfixed(0.6232)),
(re => to_ads_sfixed(0.3618) , im => to_ads_sfixed(0.6258)),
(re => to_ads_sfixed(0.3564) , im => to_ads_sfixed(0.6284)),
(re => to_ads_sfixed(0.351) , im => to_ads_sfixed(0.631)),
(re => to_ads_sfixed(0.3456) , im => to_ads_sfixed(0.6336)),
(re => to_ads_sfixed(0.3402) , im => to_ads_sfixed(0.6362)),
(re => to_ads_sfixed(0.3348) , im => to_ads_sfixed(0.6388)),
(re => to_ads_sfixed(0.3294) , im => to_ads_sfixed(0.6414)),
(re => to_ads_sfixed(0.324) , im => to_ads_sfixed(0.644)),
(re => to_ads_sfixed(0.3186) , im => to_ads_sfixed(0.6466)),
(re => to_ads_sfixed(0.3132) , im => to_ads_sfixed(0.6492)),
(re => to_ads_sfixed(0.3078) , im => to_ads_sfixed(0.6518)),
(re => to_ads_sfixed(0.3024) , im => to_ads_sfixed(0.6544)),
(re => to_ads_sfixed(0.297) , im => to_ads_sfixed(0.657)),
(re => to_ads_sfixed(0.2916) , im => to_ads_sfixed(0.6596)),
(re => to_ads_sfixed(0.2862) , im => to_ads_sfixed(0.6622)),
(re => to_ads_sfixed(0.2808) , im => to_ads_sfixed(0.6648)),
(re => to_ads_sfixed(0.2754) , im => to_ads_sfixed(0.6674)),
(re => to_ads_sfixed(0.27) , im => to_ads_sfixed(0.67)),
(re => to_ads_sfixed(0.2646) , im => to_ads_sfixed(0.6726)),
(re => to_ads_sfixed(0.2592) , im => to_ads_sfixed(0.6752)),
(re => to_ads_sfixed(0.2538) , im => to_ads_sfixed(0.6778)),
(re => to_ads_sfixed(0.2484) , im => to_ads_sfixed(0.6804)),
(re => to_ads_sfixed(0.243) , im => to_ads_sfixed(0.683)),
(re => to_ads_sfixed(0.2376) , im => to_ads_sfixed(0.6856)),
(re => to_ads_sfixed(0.2322) , im => to_ads_sfixed(0.6882)),
(re => to_ads_sfixed(0.2268) , im => to_ads_sfixed(0.6908)),
(re => to_ads_sfixed(0.2214) , im => to_ads_sfixed(0.6934)),
(re => to_ads_sfixed(0.216) , im => to_ads_sfixed(0.696)),
(re => to_ads_sfixed(0.2106) , im => to_ads_sfixed(0.6986)),
(re => to_ads_sfixed(0.2052) , im => to_ads_sfixed(0.7012)),
(re => to_ads_sfixed(0.1998) , im => to_ads_sfixed(0.7038)),
(re => to_ads_sfixed(0.1944) , im => to_ads_sfixed(0.7064)),
(re => to_ads_sfixed(0.189) , im => to_ads_sfixed(0.709)),
(re => to_ads_sfixed(0.1836) , im => to_ads_sfixed(0.7116)),
(re => to_ads_sfixed(0.1782) , im => to_ads_sfixed(0.7142)),
(re => to_ads_sfixed(0.1728) , im => to_ads_sfixed(0.7168)),
(re => to_ads_sfixed(0.1674) , im => to_ads_sfixed(0.7194)),
(re => to_ads_sfixed(0.162) , im => to_ads_sfixed(0.722)),
(re => to_ads_sfixed(0.1566) , im => to_ads_sfixed(0.7246)),
(re => to_ads_sfixed(0.1512) , im => to_ads_sfixed(0.7272)),
(re => to_ads_sfixed(0.1458) , im => to_ads_sfixed(0.7298)),
(re => to_ads_sfixed(0.1404) , im => to_ads_sfixed(0.7324)),
(re => to_ads_sfixed(0.135) , im => to_ads_sfixed(0.735)),
(re => to_ads_sfixed(0.1296) , im => to_ads_sfixed(0.7376)),
(re => to_ads_sfixed(0.1242) , im => to_ads_sfixed(0.7402)),
(re => to_ads_sfixed(0.1188) , im => to_ads_sfixed(0.7428)),
(re => to_ads_sfixed(0.1134) , im => to_ads_sfixed(0.7454)),
(re => to_ads_sfixed(0.108) , im => to_ads_sfixed(0.748)),
(re => to_ads_sfixed(0.1026) , im => to_ads_sfixed(0.7506)),
(re => to_ads_sfixed(0.0972) , im => to_ads_sfixed(0.7532)),
(re => to_ads_sfixed(0.0918) , im => to_ads_sfixed(0.7558)),
(re => to_ads_sfixed(0.0864) , im => to_ads_sfixed(0.7584)),
(re => to_ads_sfixed(0.081) , im => to_ads_sfixed(0.761)),
(re => to_ads_sfixed(0.0756) , im => to_ads_sfixed(0.7636)),
(re => to_ads_sfixed(0.0702) , im => to_ads_sfixed(0.7662)),
(re => to_ads_sfixed(0.0648) , im => to_ads_sfixed(0.7688)),
(re => to_ads_sfixed(0.0594) , im => to_ads_sfixed(0.7714)),
(re => to_ads_sfixed(0.054) , im => to_ads_sfixed(0.774)),
(re => to_ads_sfixed(0.0486) , im => to_ads_sfixed(0.7766)),
(re => to_ads_sfixed(0.0432) , im => to_ads_sfixed(0.7792)),
(re => to_ads_sfixed(0.0378) , im => to_ads_sfixed(0.7818)),
(re => to_ads_sfixed(0.0324) , im => to_ads_sfixed(0.7844)),
(re => to_ads_sfixed(0.027) , im => to_ads_sfixed(0.787)),
(re => to_ads_sfixed(0.0216) , im => to_ads_sfixed(0.7896)),
(re => to_ads_sfixed(0.0162) , im => to_ads_sfixed(0.7922)),
(re => to_ads_sfixed(0.0108) , im => to_ads_sfixed(0.7948)),
(re => to_ads_sfixed(0.0054) , im => to_ads_sfixed(0.7974)),
(re => to_ads_sfixed(0.0) , im => to_ads_sfixed(0.8)),
(re => to_ads_sfixed(-0.0054) , im => to_ads_sfixed(0.7974)),
(re => to_ads_sfixed(-0.0108) , im => to_ads_sfixed(0.7948)),
(re => to_ads_sfixed(-0.0162) , im => to_ads_sfixed(0.7922)),
(re => to_ads_sfixed(-0.0216) , im => to_ads_sfixed(0.7896)),
(re => to_ads_sfixed(-0.027) , im => to_ads_sfixed(0.787)),
(re => to_ads_sfixed(-0.0324) , im => to_ads_sfixed(0.7844)),
(re => to_ads_sfixed(-0.0378) , im => to_ads_sfixed(0.7818)),
(re => to_ads_sfixed(-0.0432) , im => to_ads_sfixed(0.7792)),
(re => to_ads_sfixed(-0.0486) , im => to_ads_sfixed(0.7766)),
(re => to_ads_sfixed(-0.054) , im => to_ads_sfixed(0.774)),
(re => to_ads_sfixed(-0.0594) , im => to_ads_sfixed(0.7714)),
(re => to_ads_sfixed(-0.0648) , im => to_ads_sfixed(0.7688)),
(re => to_ads_sfixed(-0.0702) , im => to_ads_sfixed(0.7662)),
(re => to_ads_sfixed(-0.0756) , im => to_ads_sfixed(0.7636)),
(re => to_ads_sfixed(-0.081) , im => to_ads_sfixed(0.761)),
(re => to_ads_sfixed(-0.0864) , im => to_ads_sfixed(0.7584)),
(re => to_ads_sfixed(-0.0918) , im => to_ads_sfixed(0.7558)),
(re => to_ads_sfixed(-0.0972) , im => to_ads_sfixed(0.7532)),
(re => to_ads_sfixed(-0.1026) , im => to_ads_sfixed(0.7506)),
(re => to_ads_sfixed(-0.108) , im => to_ads_sfixed(0.748)),
(re => to_ads_sfixed(-0.1134) , im => to_ads_sfixed(0.7454)),
(re => to_ads_sfixed(-0.1188) , im => to_ads_sfixed(0.7428)),
(re => to_ads_sfixed(-0.1242) , im => to_ads_sfixed(0.7402)),
(re => to_ads_sfixed(-0.1296) , im => to_ads_sfixed(0.7376)),
(re => to_ads_sfixed(-0.135) , im => to_ads_sfixed(0.735)),
(re => to_ads_sfixed(-0.1404) , im => to_ads_sfixed(0.7324)),
(re => to_ads_sfixed(-0.1458) , im => to_ads_sfixed(0.7298)),
(re => to_ads_sfixed(-0.1512) , im => to_ads_sfixed(0.7272)),
(re => to_ads_sfixed(-0.1566) , im => to_ads_sfixed(0.7246)),
(re => to_ads_sfixed(-0.162) , im => to_ads_sfixed(0.722)),
(re => to_ads_sfixed(-0.1674) , im => to_ads_sfixed(0.7194)),
(re => to_ads_sfixed(-0.1728) , im => to_ads_sfixed(0.7168)),
(re => to_ads_sfixed(-0.1782) , im => to_ads_sfixed(0.7142)),
(re => to_ads_sfixed(-0.1836) , im => to_ads_sfixed(0.7116)),
(re => to_ads_sfixed(-0.189) , im => to_ads_sfixed(0.709)),
(re => to_ads_sfixed(-0.1944) , im => to_ads_sfixed(0.7064)),
(re => to_ads_sfixed(-0.1998) , im => to_ads_sfixed(0.7038)),
(re => to_ads_sfixed(-0.2052) , im => to_ads_sfixed(0.7012)),
(re => to_ads_sfixed(-0.2106) , im => to_ads_sfixed(0.6986)),
(re => to_ads_sfixed(-0.216) , im => to_ads_sfixed(0.696)),
(re => to_ads_sfixed(-0.2214) , im => to_ads_sfixed(0.6934)),
(re => to_ads_sfixed(-0.2268) , im => to_ads_sfixed(0.6908)),
(re => to_ads_sfixed(-0.2322) , im => to_ads_sfixed(0.6882)),
(re => to_ads_sfixed(-0.2376) , im => to_ads_sfixed(0.6856)),
(re => to_ads_sfixed(-0.243) , im => to_ads_sfixed(0.683)),
(re => to_ads_sfixed(-0.2484) , im => to_ads_sfixed(0.6804)),
(re => to_ads_sfixed(-0.2538) , im => to_ads_sfixed(0.6778)),
(re => to_ads_sfixed(-0.2592) , im => to_ads_sfixed(0.6752)),
(re => to_ads_sfixed(-0.2646) , im => to_ads_sfixed(0.6726)),
(re => to_ads_sfixed(-0.27) , im => to_ads_sfixed(0.67)),
(re => to_ads_sfixed(-0.2754) , im => to_ads_sfixed(0.6674)),
(re => to_ads_sfixed(-0.2808) , im => to_ads_sfixed(0.6648)),
(re => to_ads_sfixed(-0.2862) , im => to_ads_sfixed(0.6622)),
(re => to_ads_sfixed(-0.2916) , im => to_ads_sfixed(0.6596)),
(re => to_ads_sfixed(-0.297) , im => to_ads_sfixed(0.657)),
(re => to_ads_sfixed(-0.3024) , im => to_ads_sfixed(0.6544)),
(re => to_ads_sfixed(-0.3078) , im => to_ads_sfixed(0.6518)),
(re => to_ads_sfixed(-0.3132) , im => to_ads_sfixed(0.6492)),
(re => to_ads_sfixed(-0.3186) , im => to_ads_sfixed(0.6466)),
(re => to_ads_sfixed(-0.324) , im => to_ads_sfixed(0.644)),
(re => to_ads_sfixed(-0.3294) , im => to_ads_sfixed(0.6414)),
(re => to_ads_sfixed(-0.3348) , im => to_ads_sfixed(0.6388)),
(re => to_ads_sfixed(-0.3402) , im => to_ads_sfixed(0.6362)),
(re => to_ads_sfixed(-0.3456) , im => to_ads_sfixed(0.6336)),
(re => to_ads_sfixed(-0.351) , im => to_ads_sfixed(0.631)),
(re => to_ads_sfixed(-0.3564) , im => to_ads_sfixed(0.6284)),
(re => to_ads_sfixed(-0.3618) , im => to_ads_sfixed(0.6258)),
(re => to_ads_sfixed(-0.3672) , im => to_ads_sfixed(0.6232)),
(re => to_ads_sfixed(-0.3726) , im => to_ads_sfixed(0.6206)),
(re => to_ads_sfixed(-0.378) , im => to_ads_sfixed(0.618)),
(re => to_ads_sfixed(-0.3834) , im => to_ads_sfixed(0.6154)),
(re => to_ads_sfixed(-0.3888) , im => to_ads_sfixed(0.6128)),
(re => to_ads_sfixed(-0.3942) , im => to_ads_sfixed(0.6102)),
(re => to_ads_sfixed(-0.3996) , im => to_ads_sfixed(0.6076)),
(re => to_ads_sfixed(-0.405) , im => to_ads_sfixed(0.605)),
(re => to_ads_sfixed(-0.4104) , im => to_ads_sfixed(0.6024)),
(re => to_ads_sfixed(-0.4158) , im => to_ads_sfixed(0.5998)),
(re => to_ads_sfixed(-0.4212) , im => to_ads_sfixed(0.5972)),
(re => to_ads_sfixed(-0.4266) , im => to_ads_sfixed(0.5946)),
(re => to_ads_sfixed(-0.432) , im => to_ads_sfixed(0.592)),
(re => to_ads_sfixed(-0.4374) , im => to_ads_sfixed(0.5894)),
(re => to_ads_sfixed(-0.4428) , im => to_ads_sfixed(0.5868)),
(re => to_ads_sfixed(-0.4482) , im => to_ads_sfixed(0.5842)),
(re => to_ads_sfixed(-0.4536) , im => to_ads_sfixed(0.5816)),
(re => to_ads_sfixed(-0.459) , im => to_ads_sfixed(0.579)),
(re => to_ads_sfixed(-0.4644) , im => to_ads_sfixed(0.5764)),
(re => to_ads_sfixed(-0.4698) , im => to_ads_sfixed(0.5738)),
(re => to_ads_sfixed(-0.4752) , im => to_ads_sfixed(0.5712)),
(re => to_ads_sfixed(-0.4806) , im => to_ads_sfixed(0.5686)),
(re => to_ads_sfixed(-0.486) , im => to_ads_sfixed(0.566)),
(re => to_ads_sfixed(-0.4914) , im => to_ads_sfixed(0.5634)),
(re => to_ads_sfixed(-0.4968) , im => to_ads_sfixed(0.5608)),
(re => to_ads_sfixed(-0.5022) , im => to_ads_sfixed(0.5582)),
(re => to_ads_sfixed(-0.5076) , im => to_ads_sfixed(0.5556)),
(re => to_ads_sfixed(-0.513) , im => to_ads_sfixed(0.553)),
(re => to_ads_sfixed(-0.5184) , im => to_ads_sfixed(0.5504)),
(re => to_ads_sfixed(-0.5238) , im => to_ads_sfixed(0.5478)),
(re => to_ads_sfixed(-0.5292) , im => to_ads_sfixed(0.5452)),
(re => to_ads_sfixed(-0.5346) , im => to_ads_sfixed(0.5426)),
(re => to_ads_sfixed(-0.54) , im => to_ads_sfixed(0.54)),
(re => to_ads_sfixed(-0.5362) , im => to_ads_sfixed(0.545005)),
(re => to_ads_sfixed(-0.5324) , im => to_ads_sfixed(0.55001)),
(re => to_ads_sfixed(-0.5286) , im => to_ads_sfixed(0.555015)),
(re => to_ads_sfixed(-0.5248) , im => to_ads_sfixed(0.56002)),
(re => to_ads_sfixed(-0.521) , im => to_ads_sfixed(0.565025)),
(re => to_ads_sfixed(-0.5172) , im => to_ads_sfixed(0.57003)),
(re => to_ads_sfixed(-0.5134) , im => to_ads_sfixed(0.575035)),
(re => to_ads_sfixed(-0.5096) , im => to_ads_sfixed(0.58004)),
(re => to_ads_sfixed(-0.5058) , im => to_ads_sfixed(0.585045)),
(re => to_ads_sfixed(-0.502) , im => to_ads_sfixed(0.59005)),
(re => to_ads_sfixed(-0.4982) , im => to_ads_sfixed(0.595055)),
(re => to_ads_sfixed(-0.4944) , im => to_ads_sfixed(0.60006)),
(re => to_ads_sfixed(-0.4906) , im => to_ads_sfixed(0.605065)),
(re => to_ads_sfixed(-0.4868) , im => to_ads_sfixed(0.61007)),
(re => to_ads_sfixed(-0.483) , im => to_ads_sfixed(0.615075)),
(re => to_ads_sfixed(-0.4792) , im => to_ads_sfixed(0.62008)),
(re => to_ads_sfixed(-0.4754) , im => to_ads_sfixed(0.625085)),
(re => to_ads_sfixed(-0.4716) , im => to_ads_sfixed(0.63009)),
(re => to_ads_sfixed(-0.4678) , im => to_ads_sfixed(0.635095)),
(re => to_ads_sfixed(-0.464) , im => to_ads_sfixed(0.6401)),
(re => to_ads_sfixed(-0.4602) , im => to_ads_sfixed(0.645105)),
(re => to_ads_sfixed(-0.4564) , im => to_ads_sfixed(0.65011)),
(re => to_ads_sfixed(-0.4526) , im => to_ads_sfixed(0.655115)),
(re => to_ads_sfixed(-0.4488) , im => to_ads_sfixed(0.66012)),
(re => to_ads_sfixed(-0.445) , im => to_ads_sfixed(0.665125)),
(re => to_ads_sfixed(-0.4412) , im => to_ads_sfixed(0.67013)),
(re => to_ads_sfixed(-0.4374) , im => to_ads_sfixed(0.675135)),
(re => to_ads_sfixed(-0.4336) , im => to_ads_sfixed(0.68014)),
(re => to_ads_sfixed(-0.4298) , im => to_ads_sfixed(0.685145)),
(re => to_ads_sfixed(-0.426) , im => to_ads_sfixed(0.69015)),
(re => to_ads_sfixed(-0.4222) , im => to_ads_sfixed(0.695155)),
(re => to_ads_sfixed(-0.4184) , im => to_ads_sfixed(0.70016)),
(re => to_ads_sfixed(-0.4146) , im => to_ads_sfixed(0.705165)),
(re => to_ads_sfixed(-0.4108) , im => to_ads_sfixed(0.71017)),
(re => to_ads_sfixed(-0.407) , im => to_ads_sfixed(0.715175)),
(re => to_ads_sfixed(-0.4032) , im => to_ads_sfixed(0.72018)),
(re => to_ads_sfixed(-0.3994) , im => to_ads_sfixed(0.725185)),
(re => to_ads_sfixed(-0.3956) , im => to_ads_sfixed(0.73019)),
(re => to_ads_sfixed(-0.3918) , im => to_ads_sfixed(0.735195)),
(re => to_ads_sfixed(-0.388) , im => to_ads_sfixed(0.7402)),
(re => to_ads_sfixed(-0.3842) , im => to_ads_sfixed(0.745205)),
(re => to_ads_sfixed(-0.3804) , im => to_ads_sfixed(0.75021)),
(re => to_ads_sfixed(-0.3766) , im => to_ads_sfixed(0.755215)),
(re => to_ads_sfixed(-0.3728) , im => to_ads_sfixed(0.76022)),
(re => to_ads_sfixed(-0.369) , im => to_ads_sfixed(0.765225)),
(re => to_ads_sfixed(-0.3652) , im => to_ads_sfixed(0.77023)),
(re => to_ads_sfixed(-0.3614) , im => to_ads_sfixed(0.775235)),
(re => to_ads_sfixed(-0.3576) , im => to_ads_sfixed(0.78024)),
(re => to_ads_sfixed(-0.3538) , im => to_ads_sfixed(0.785245)),
(re => to_ads_sfixed(-0.35) , im => to_ads_sfixed(0.79025)),
(re => to_ads_sfixed(-0.3462) , im => to_ads_sfixed(0.795255)),
(re => to_ads_sfixed(-0.3424) , im => to_ads_sfixed(0.80026)),
(re => to_ads_sfixed(-0.3386) , im => to_ads_sfixed(0.805265)),
(re => to_ads_sfixed(-0.3348) , im => to_ads_sfixed(0.81027)),
(re => to_ads_sfixed(-0.331) , im => to_ads_sfixed(0.815275)),
(re => to_ads_sfixed(-0.3272) , im => to_ads_sfixed(0.82028)),
(re => to_ads_sfixed(-0.3234) , im => to_ads_sfixed(0.825285)),
(re => to_ads_sfixed(-0.3196) , im => to_ads_sfixed(0.83029)),
(re => to_ads_sfixed(-0.3158) , im => to_ads_sfixed(0.835295)),
(re => to_ads_sfixed(-0.312) , im => to_ads_sfixed(0.8403)),
(re => to_ads_sfixed(-0.3082) , im => to_ads_sfixed(0.845305)),
(re => to_ads_sfixed(-0.3044) , im => to_ads_sfixed(0.85031)),
(re => to_ads_sfixed(-0.3006) , im => to_ads_sfixed(0.855315)),
(re => to_ads_sfixed(-0.2968) , im => to_ads_sfixed(0.86032)),
(re => to_ads_sfixed(-0.293) , im => to_ads_sfixed(0.865325)),
(re => to_ads_sfixed(-0.2892) , im => to_ads_sfixed(0.87033)),
(re => to_ads_sfixed(-0.2854) , im => to_ads_sfixed(0.875335)),
(re => to_ads_sfixed(-0.2816) , im => to_ads_sfixed(0.88034)),
(re => to_ads_sfixed(-0.2778) , im => to_ads_sfixed(0.885345)),
(re => to_ads_sfixed(-0.274) , im => to_ads_sfixed(0.89035)),
(re => to_ads_sfixed(-0.2702) , im => to_ads_sfixed(0.895355)),
(re => to_ads_sfixed(-0.2664) , im => to_ads_sfixed(0.90036)),
(re => to_ads_sfixed(-0.2626) , im => to_ads_sfixed(0.905365)),
(re => to_ads_sfixed(-0.2588) , im => to_ads_sfixed(0.91037)),
(re => to_ads_sfixed(-0.255) , im => to_ads_sfixed(0.915375)),
(re => to_ads_sfixed(-0.2512) , im => to_ads_sfixed(0.92038)),
(re => to_ads_sfixed(-0.2474) , im => to_ads_sfixed(0.925385)),
(re => to_ads_sfixed(-0.2436) , im => to_ads_sfixed(0.93039)),
(re => to_ads_sfixed(-0.2398) , im => to_ads_sfixed(0.935395)),
(re => to_ads_sfixed(-0.236) , im => to_ads_sfixed(0.9404)),
(re => to_ads_sfixed(-0.2322) , im => to_ads_sfixed(0.945405)),
(re => to_ads_sfixed(-0.2284) , im => to_ads_sfixed(0.95041)),
(re => to_ads_sfixed(-0.2246) , im => to_ads_sfixed(0.955415)),
(re => to_ads_sfixed(-0.2208) , im => to_ads_sfixed(0.96042)),
(re => to_ads_sfixed(-0.217) , im => to_ads_sfixed(0.965425)),
(re => to_ads_sfixed(-0.2132) , im => to_ads_sfixed(0.97043)),
(re => to_ads_sfixed(-0.2094) , im => to_ads_sfixed(0.975435)),
(re => to_ads_sfixed(-0.2056) , im => to_ads_sfixed(0.98044)),
(re => to_ads_sfixed(-0.2018) , im => to_ads_sfixed(0.985445)),
(re => to_ads_sfixed(-0.198) , im => to_ads_sfixed(0.99045)),
(re => to_ads_sfixed(-0.1942) , im => to_ads_sfixed(0.995455)),
(re => to_ads_sfixed(-0.1904) , im => to_ads_sfixed(1.00046)),
(re => to_ads_sfixed(-0.1866) , im => to_ads_sfixed(1.005465)),
(re => to_ads_sfixed(-0.1828) , im => to_ads_sfixed(1.01047)),
(re => to_ads_sfixed(-0.179) , im => to_ads_sfixed(1.015475)),
(re => to_ads_sfixed(-0.1752) , im => to_ads_sfixed(1.02048)),
(re => to_ads_sfixed(-0.1714) , im => to_ads_sfixed(1.025485)),
(re => to_ads_sfixed(-0.1676) , im => to_ads_sfixed(1.03049)),
(re => to_ads_sfixed(-0.1638) , im => to_ads_sfixed(1.035495))); 	
		
end package mandlebrot_pkg;

package body mandlebrot_pkg is

end package body mandlebrot_pkg;