* ring_oscillator_2

.include nand.cir
.include inverter.cir

.subckt ring_oscillator_2 in out vdd vss
x0 in out s1 vdd vss nand
x1 s1 s2 vdd vss inverter tplv=6.103918639686384e-08 tpwv=2.0669282684218656e-07 tnln=6.895137477075377e-08 tnwn=1.1101954929680408e-07 tpotv=2.036899030671505e-09 tnotv=1.9510379806218446e-09 inverter
x2 s2 s3 vdd vss inverter tplv=6.964055514470665e-08 tpwv=2.214073622689235e-07 tnln=6.04844626492672e-08 tnwn=1.3607719133329308e-07 tpotv=2.099848689315428e-09 tnotv=1.9599025102501486e-09 inverter
x3 s3 s4 vdd vss inverter tplv=6.426775385339483e-08 tpwv=2.122985230590509e-07 tnln=6.311342074510594e-08 tnwn=1.1587854200384855e-07 tpotv=2.0322267982508322e-09 tnotv=1.6825744230726994e-09 inverter
x4 s4 s5 vdd vss inverter tplv=6.431045525761368e-08 tpwv=2.2075475937266273e-07 tnln=7.546471410361156e-08 tnwn=1.3416468459910032e-07 tpotv=1.980773387656511e-09 tnotv=1.884685581795874e-09 inverter
x5 s5 s6 vdd vss inverter tplv=6.479920665527815e-08 tpwv=2.0405630405071017e-07 tnln=7.383430569021665e-08 tnwn=1.2720354504535223e-07 tpotv=1.927465325180225e-09 tnotv=1.9514455434045765e-09 inverter
x6 s6 s7 vdd vss inverter tplv=6.383495759392275e-08 tpwv=2.0487042958726507e-07 tnln=6.603951373439844e-08 tnwn=1.34828001267717e-07 tpotv=1.8728491069906075e-09 tnotv=1.935916288468687e-09 inverter
x7 s7 s8 vdd vss inverter tplv=6.922506734353715e-08 tpwv=2.159661595865519e-07 tnln=5.614708144410589e-08 tnwn=1.3941842881834413e-07 tpotv=1.9647819082579667e-09 tnotv=1.775138724181785e-09 inverter
x8 s8 s9 vdd vss inverter tplv=6.245414319193241e-08 tpwv=2.1432590826448558e-07 tnln=6.473404995911516e-08 tnwn=1.0404314136541422e-07 tpotv=1.841441659872306e-09 tnotv=1.8901899858408567e-09 inverter
x9 s9 s10 vdd vss inverter tplv=7.422986553743817e-08 tpwv=2.0018645223173968e-07 tnln=6.079984650700142e-08 tnwn=1.3325353209436207e-07 tpotv=2.017056213001008e-09 tnotv=1.8965412464492107e-09 inverter
x10 s10 s11 vdd vss inverter tplv=6.083823681978555e-08 tpwv=2.1759365058933406e-07 tnln=6.145361693849844e-08 tnwn=1.2334520693865735e-07 tpotv=1.8023006377278987e-09 tnotv=1.9213930934993855e-09 inverter
x11 s11 s12 vdd vss inverter tplv=6.455634557781755e-08 tpwv=1.9838873717139663e-07 tnln=6.329637995005493e-08 tnwn=1.3680330563865652e-07 tpotv=1.959157299955536e-09 tnotv=1.7412216022753487e-09 inverter
x12 s12 out vdd vss inverter tplv=6.58853867691965e-08 tpwv=2.0577151649904824e-07 tnln=6.06129420567889e-08 tnwn=1.1605829319668854e-07 tpotv=1.9690920320235018e-09 tnotv=1.710452967705821e-09 inverter
.ends ring_oscillator_2